// Testbench

`timescale 1ns / 1ps

module tb_Top;

    reg clk;
    reg reset;
    reg signed [7:0] A; 
    reg signed [7:0] B;
    wire signed [15:0] Output;

    Top uut (
        .clk(clk), 
        .reset(reset), 
        .A(A), 
        .B(B), 
        .Output(Output)
    );

    initial begin
        clk = 0;
        forever #5 clk = ~clk; 
    end

    initial begin

        $monitor("Time=%0t | Input: %d * %d | Output=%d ", 
                 $time, A, B, Output);

  
        reset = 1; A = 0; B = 0;
        #100;  // wait for global reset (100ns)
        #15;
        reset = 0;
        #1;

        // ------------------------------------------------------------
        // Test Case 1: Positive * Positive (4 * 5 = 20)
        // ------------------------------------------------------------
        A = 4; B = 5;
        #20; // Wait for pipeline

        // ------------------------------------------------------------
        // Test Case 2: Positive * Negative (10 * -2 = -20)
        // ------------------------------------------------------------
        A = 10; B = -2;
        #20;

        // ------------------------------------------------------------
        // Test Case 3: Negative * Positive (-5 * 5 = -25)
        // ------------------------------------------------------------
        A = -5; B = 5;
        #20;

        // ------------------------------------------------------------
        // Test Case 4: Negative * Negative (-10 * -10 = 100)
        // ------------------------------------------------------------
        A = -10; B = -10;
        #20;

        // ------------------------------------------------------------
        // Test Case 5: Max Boundary Test (127 * 127 = 16129)
        // ------------------------------------------------------------
        A = 127; B = 127;
        #20;

        // ------------------------------------------------------------
        // Test Case 6: Min Boundary Test (-128 * 1 = -128)
        // ------------------------------------------------------------
        A = -128; B = 1;
        #50;

        $finish;
    end

endmodule