VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Top
  CLASS BLOCK ;
  FOREIGN Top ;
  ORIGIN 0.000 0.000 ;
  SIZE 94.785 BY 105.505 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 5.610 101.505 5.890 105.505 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 11.130 101.505 11.410 105.505 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 16.650 101.505 16.930 105.505 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 22.170 101.505 22.450 105.505 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 27.690 101.505 27.970 105.505 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 33.210 101.505 33.490 105.505 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 101.505 39.010 105.505 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 44.250 101.505 44.530 105.505 ;
    END
  END A[7]
  PIN B[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 49.770 101.505 50.050 105.505 ;
    END
  END B[0]
  PIN B[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 55.290 101.505 55.570 105.505 ;
    END
  END B[1]
  PIN B[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 60.810 101.505 61.090 105.505 ;
    END
  END B[2]
  PIN B[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 66.330 101.505 66.610 105.505 ;
    END
  END B[3]
  PIN B[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 71.850 101.505 72.130 105.505 ;
    END
  END B[4]
  PIN B[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 77.370 101.505 77.650 105.505 ;
    END
  END B[5]
  PIN B[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 82.890 101.505 83.170 105.505 ;
    END
  END B[6]
  PIN B[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 88.410 101.505 88.690 105.505 ;
    END
  END B[7]
  PIN Output[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END Output[0]
  PIN Output[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END Output[10]
  PIN Output[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END Output[11]
  PIN Output[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END Output[12]
  PIN Output[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END Output[13]
  PIN Output[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END Output[14]
  PIN Output[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END Output[15]
  PIN Output[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END Output[1]
  PIN Output[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END Output[2]
  PIN Output[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END Output[3]
  PIN Output[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END Output[4]
  PIN Output[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END Output[5]
  PIN Output[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END Output[6]
  PIN Output[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END Output[7]
  PIN Output[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END Output[8]
  PIN Output[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.340600 ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END Output[9]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 13.220 10.640 15.220 92.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 43.220 10.640 45.220 92.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.220 10.640 75.220 92.720 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 18.580 89.480 20.580 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 48.580 89.480 50.580 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 78.580 89.480 80.580 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.520 10.640 11.520 92.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 39.520 10.640 41.520 92.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 69.520 10.640 71.520 92.720 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 14.880 89.480 16.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 44.880 89.480 46.880 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 74.880 89.480 76.880 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 90.785 51.720 94.785 52.320 ;
    END
  END clk
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END reset
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 89.430 92.565 ;
      LAYER li1 ;
        RECT 5.520 10.795 89.240 92.565 ;
      LAYER met1 ;
        RECT 4.210 10.640 89.240 92.720 ;
      LAYER met2 ;
        RECT 4.230 101.225 5.330 101.730 ;
        RECT 6.170 101.225 10.850 101.730 ;
        RECT 11.690 101.225 16.370 101.730 ;
        RECT 17.210 101.225 21.890 101.730 ;
        RECT 22.730 101.225 27.410 101.730 ;
        RECT 28.250 101.225 32.930 101.730 ;
        RECT 33.770 101.225 38.450 101.730 ;
        RECT 39.290 101.225 43.970 101.730 ;
        RECT 44.810 101.225 49.490 101.730 ;
        RECT 50.330 101.225 55.010 101.730 ;
        RECT 55.850 101.225 60.530 101.730 ;
        RECT 61.370 101.225 66.050 101.730 ;
        RECT 66.890 101.225 71.570 101.730 ;
        RECT 72.410 101.225 77.090 101.730 ;
        RECT 77.930 101.225 82.610 101.730 ;
        RECT 83.450 101.225 88.130 101.730 ;
        RECT 4.230 4.280 88.680 101.225 ;
        RECT 4.230 4.000 46.730 4.280 ;
        RECT 47.570 4.000 88.680 4.280 ;
      LAYER met3 ;
        RECT 4.400 92.120 90.785 92.985 ;
        RECT 3.990 88.080 90.785 92.120 ;
        RECT 4.400 86.680 90.785 88.080 ;
        RECT 3.990 82.640 90.785 86.680 ;
        RECT 4.400 81.240 90.785 82.640 ;
        RECT 3.990 77.200 90.785 81.240 ;
        RECT 4.400 75.800 90.785 77.200 ;
        RECT 3.990 71.760 90.785 75.800 ;
        RECT 4.400 70.360 90.785 71.760 ;
        RECT 3.990 66.320 90.785 70.360 ;
        RECT 4.400 64.920 90.785 66.320 ;
        RECT 3.990 60.880 90.785 64.920 ;
        RECT 4.400 59.480 90.785 60.880 ;
        RECT 3.990 55.440 90.785 59.480 ;
        RECT 4.400 54.040 90.785 55.440 ;
        RECT 3.990 52.720 90.785 54.040 ;
        RECT 3.990 51.320 90.385 52.720 ;
        RECT 3.990 50.000 90.785 51.320 ;
        RECT 4.400 48.600 90.785 50.000 ;
        RECT 3.990 44.560 90.785 48.600 ;
        RECT 4.400 43.160 90.785 44.560 ;
        RECT 3.990 39.120 90.785 43.160 ;
        RECT 4.400 37.720 90.785 39.120 ;
        RECT 3.990 33.680 90.785 37.720 ;
        RECT 4.400 32.280 90.785 33.680 ;
        RECT 3.990 28.240 90.785 32.280 ;
        RECT 4.400 26.840 90.785 28.240 ;
        RECT 3.990 22.800 90.785 26.840 ;
        RECT 4.400 21.400 90.785 22.800 ;
        RECT 3.990 17.360 90.785 21.400 ;
        RECT 4.400 15.960 90.785 17.360 ;
        RECT 3.990 11.920 90.785 15.960 ;
        RECT 4.400 10.715 90.785 11.920 ;
      LAYER met4 ;
        RECT 62.855 32.135 69.120 90.265 ;
        RECT 71.920 32.135 72.385 90.265 ;
  END
END Top
END LIBRARY

