module Top (clk,
    reset,
    A,
    B,
    Output);
 input clk;
 input reset;
 input [7:0] A;
 input [7:0] B;
 output [15:0] Output;

 wire \A_ff[0] ;
 wire \A_ff[1] ;
 wire \A_ff[2] ;
 wire \A_ff[3] ;
 wire \A_ff[4] ;
 wire \A_ff[5] ;
 wire \A_ff[6] ;
 wire \A_ff[7] ;
 wire \Adder.cla_16_bit.Sum[0] ;
 wire \Adder.cla_16_bit.Sum[10] ;
 wire \Adder.cla_16_bit.Sum[11] ;
 wire \Adder.cla_16_bit.Sum[12] ;
 wire \Adder.cla_16_bit.Sum[13] ;
 wire \Adder.cla_16_bit.Sum[14] ;
 wire \Adder.cla_16_bit.Sum[15] ;
 wire \Adder.cla_16_bit.Sum[1] ;
 wire \Adder.cla_16_bit.Sum[2] ;
 wire \Adder.cla_16_bit.Sum[3] ;
 wire \Adder.cla_16_bit.Sum[4] ;
 wire \Adder.cla_16_bit.Sum[5] ;
 wire \Adder.cla_16_bit.Sum[6] ;
 wire \Adder.cla_16_bit.Sum[7] ;
 wire \Adder.cla_16_bit.Sum[8] ;
 wire \Adder.cla_16_bit.Sum[9] ;
 wire \B_ff[0] ;
 wire \B_ff[1] ;
 wire \B_ff[2] ;
 wire \B_ff[3] ;
 wire \B_ff[4] ;
 wire \B_ff[5] ;
 wire \B_ff[6] ;
 wire \B_ff[7] ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 sky130_fd_sc_hd__inv_2 _313_ (.A(\A_ff[0] ),
    .Y(_283_));
 sky130_fd_sc_hd__inv_2 _314_ (.A(\A_ff[2] ),
    .Y(_284_));
 sky130_fd_sc_hd__inv_2 _315_ (.A(\A_ff[4] ),
    .Y(_285_));
 sky130_fd_sc_hd__inv_2 _316_ (.A(\A_ff[6] ),
    .Y(_286_));
 sky130_fd_sc_hd__inv_2 _317_ (.A(\A_ff[7] ),
    .Y(_287_));
 sky130_fd_sc_hd__inv_2 _318_ (.A(net17),
    .Y(_000_));
 sky130_fd_sc_hd__and2_1 _319_ (.A(\B_ff[0] ),
    .B(\A_ff[0] ),
    .X(\Adder.cla_16_bit.Sum[0] ));
 sky130_fd_sc_hd__nand2_1 _320_ (.A(\B_ff[0] ),
    .B(\A_ff[1] ),
    .Y(_288_));
 sky130_fd_sc_hd__nand2_1 _321_ (.A(\B_ff[1] ),
    .B(\A_ff[0] ),
    .Y(_289_));
 sky130_fd_sc_hd__xor2_1 _322_ (.A(_288_),
    .B(_289_),
    .X(\Adder.cla_16_bit.Sum[1] ));
 sky130_fd_sc_hd__and2_1 _323_ (.A(\B_ff[0] ),
    .B(\B_ff[1] ),
    .X(_290_));
 sky130_fd_sc_hd__nand2_1 _324_ (.A(\B_ff[0] ),
    .B(\B_ff[1] ),
    .Y(_291_));
 sky130_fd_sc_hd__nand2b_2 _325_ (.A_N(\B_ff[0] ),
    .B(\B_ff[1] ),
    .Y(_292_));
 sky130_fd_sc_hd__and2b_1 _326_ (.A_N(\B_ff[1] ),
    .B(\B_ff[0] ),
    .X(_293_));
 sky130_fd_sc_hd__nand2b_1 _327_ (.A_N(\B_ff[1] ),
    .B(\B_ff[0] ),
    .Y(_294_));
 sky130_fd_sc_hd__nand2_1 _328_ (.A(\A_ff[2] ),
    .B(_293_),
    .Y(_295_));
 sky130_fd_sc_hd__o221a_1 _329_ (.A1(\A_ff[2] ),
    .A2(_291_),
    .B1(_292_),
    .B2(\A_ff[1] ),
    .C1(_295_),
    .X(_296_));
 sky130_fd_sc_hd__and3_1 _330_ (.A(\B_ff[1] ),
    .B(_283_),
    .C(_288_),
    .X(_297_));
 sky130_fd_sc_hd__nand2_1 _331_ (.A(\B_ff[1] ),
    .B(\B_ff[2] ),
    .Y(_298_));
 sky130_fd_sc_hd__xnor2_4 _332_ (.A(\B_ff[1] ),
    .B(\B_ff[2] ),
    .Y(_299_));
 sky130_fd_sc_hd__inv_2 _333_ (.A(_299_),
    .Y(_300_));
 sky130_fd_sc_hd__a21o_1 _334_ (.A1(\A_ff[0] ),
    .A2(_300_),
    .B1(_297_),
    .X(_301_));
 sky130_fd_sc_hd__xnor2_1 _335_ (.A(_296_),
    .B(_301_),
    .Y(\Adder.cla_16_bit.Sum[2] ));
 sky130_fd_sc_hd__nand2b_1 _336_ (.A_N(_296_),
    .B(_297_),
    .Y(_302_));
 sky130_fd_sc_hd__a21boi_1 _337_ (.A1(\B_ff[1] ),
    .A2(\B_ff[2] ),
    .B1_N(\B_ff[3] ),
    .Y(_303_));
 sky130_fd_sc_hd__a21oi_1 _338_ (.A1(\A_ff[0] ),
    .A2(_300_),
    .B1(_303_),
    .Y(_304_));
 sky130_fd_sc_hd__nor3b_1 _339_ (.A(\B_ff[1] ),
    .B(\B_ff[2] ),
    .C_N(\B_ff[3] ),
    .Y(_305_));
 sky130_fd_sc_hd__or3b_1 _340_ (.A(\B_ff[1] ),
    .B(\B_ff[2] ),
    .C_N(\B_ff[3] ),
    .X(_306_));
 sky130_fd_sc_hd__a31o_1 _341_ (.A1(\A_ff[0] ),
    .A2(_296_),
    .A3(_306_),
    .B1(_304_),
    .X(_307_));
 sky130_fd_sc_hd__mux2_1 _342_ (.A0(_291_),
    .A1(_294_),
    .S(\A_ff[3] ),
    .X(_308_));
 sky130_fd_sc_hd__o21ai_2 _343_ (.A1(\A_ff[2] ),
    .A2(_292_),
    .B1(_308_),
    .Y(_309_));
 sky130_fd_sc_hd__a2bb2o_1 _344_ (.A1_N(\A_ff[1] ),
    .A2_N(_299_),
    .B1(_305_),
    .B2(_283_),
    .X(_310_));
 sky130_fd_sc_hd__o21ba_1 _345_ (.A1(\B_ff[1] ),
    .A2(\B_ff[2] ),
    .B1_N(\B_ff[3] ),
    .X(_311_));
 sky130_fd_sc_hd__o21bai_1 _346_ (.A1(\B_ff[1] ),
    .A2(\B_ff[2] ),
    .B1_N(\B_ff[3] ),
    .Y(_312_));
 sky130_fd_sc_hd__or2_2 _347_ (.A(\B_ff[3] ),
    .B(_299_),
    .X(_032_));
 sky130_fd_sc_hd__o21a_1 _348_ (.A1(\A_ff[0] ),
    .A2(_298_),
    .B1(_311_),
    .X(_033_));
 sky130_fd_sc_hd__o22a_1 _349_ (.A1(\A_ff[1] ),
    .A2(_032_),
    .B1(_033_),
    .B2(_310_),
    .X(_034_));
 sky130_fd_sc_hd__nand2_1 _350_ (.A(_309_),
    .B(_034_),
    .Y(_035_));
 sky130_fd_sc_hd__nor2_1 _351_ (.A(_309_),
    .B(_034_),
    .Y(_036_));
 sky130_fd_sc_hd__xnor2_1 _352_ (.A(_309_),
    .B(_034_),
    .Y(_037_));
 sky130_fd_sc_hd__a21oi_1 _353_ (.A1(_307_),
    .A2(_035_),
    .B1(_036_),
    .Y(_038_));
 sky130_fd_sc_hd__xor2_1 _354_ (.A(_307_),
    .B(_037_),
    .X(_039_));
 sky130_fd_sc_hd__and2b_1 _355_ (.A_N(_302_),
    .B(_039_),
    .X(_040_));
 sky130_fd_sc_hd__xnor2_1 _356_ (.A(_302_),
    .B(_039_),
    .Y(\Adder.cla_16_bit.Sum[3] ));
 sky130_fd_sc_hd__and2_1 _357_ (.A(\B_ff[3] ),
    .B(\B_ff[4] ),
    .X(_041_));
 sky130_fd_sc_hd__nand2_1 _358_ (.A(\B_ff[3] ),
    .B(\B_ff[4] ),
    .Y(_042_));
 sky130_fd_sc_hd__a21bo_1 _359_ (.A1(\B_ff[3] ),
    .A2(\B_ff[4] ),
    .B1_N(\B_ff[5] ),
    .X(_043_));
 sky130_fd_sc_hd__nor2_1 _360_ (.A(\B_ff[3] ),
    .B(\B_ff[4] ),
    .Y(_044_));
 sky130_fd_sc_hd__o21ba_1 _361_ (.A1(\B_ff[3] ),
    .A2(\B_ff[4] ),
    .B1_N(\B_ff[5] ),
    .X(_045_));
 sky130_fd_sc_hd__o21bai_2 _362_ (.A1(\B_ff[3] ),
    .A2(\B_ff[4] ),
    .B1_N(\B_ff[5] ),
    .Y(_046_));
 sky130_fd_sc_hd__nand2_1 _363_ (.A(\A_ff[0] ),
    .B(_045_),
    .Y(_047_));
 sky130_fd_sc_hd__o21ai_1 _364_ (.A1(_283_),
    .A2(_044_),
    .B1(\B_ff[5] ),
    .Y(_048_));
 sky130_fd_sc_hd__a21oi_1 _365_ (.A1(_047_),
    .A2(_048_),
    .B1(_041_),
    .Y(_049_));
 sky130_fd_sc_hd__nand3b_1 _366_ (.A_N(\B_ff[1] ),
    .B(\A_ff[4] ),
    .C(\B_ff[0] ),
    .Y(_050_));
 sky130_fd_sc_hd__o221a_1 _367_ (.A1(\A_ff[4] ),
    .A2(_291_),
    .B1(_292_),
    .B2(\A_ff[3] ),
    .C1(_050_),
    .X(_051_));
 sky130_fd_sc_hd__and3b_1 _368_ (.A_N(\A_ff[1] ),
    .B(\B_ff[2] ),
    .C(\B_ff[1] ),
    .X(_052_));
 sky130_fd_sc_hd__or4b_1 _369_ (.A(\B_ff[1] ),
    .B(\A_ff[1] ),
    .C(\B_ff[2] ),
    .D_N(\B_ff[3] ),
    .X(_053_));
 sky130_fd_sc_hd__o221ai_2 _370_ (.A1(\A_ff[2] ),
    .A2(_299_),
    .B1(_312_),
    .B2(_052_),
    .C1(_053_),
    .Y(_054_));
 sky130_fd_sc_hd__or3_1 _371_ (.A(\A_ff[2] ),
    .B(\B_ff[3] ),
    .C(_299_),
    .X(_055_));
 sky130_fd_sc_hd__nand3b_1 _372_ (.A_N(_051_),
    .B(_054_),
    .C(_055_),
    .Y(_056_));
 sky130_fd_sc_hd__a21bo_1 _373_ (.A1(_054_),
    .A2(_055_),
    .B1_N(_051_),
    .X(_057_));
 sky130_fd_sc_hd__a21oi_1 _374_ (.A1(_056_),
    .A2(_057_),
    .B1(_049_),
    .Y(_058_));
 sky130_fd_sc_hd__and3_1 _375_ (.A(_049_),
    .B(_056_),
    .C(_057_),
    .X(_059_));
 sky130_fd_sc_hd__or3_2 _376_ (.A(_043_),
    .B(_058_),
    .C(_059_),
    .X(_060_));
 sky130_fd_sc_hd__o21ai_1 _377_ (.A1(_058_),
    .A2(_059_),
    .B1(_043_),
    .Y(_061_));
 sky130_fd_sc_hd__and3_1 _378_ (.A(_038_),
    .B(_060_),
    .C(_061_),
    .X(_062_));
 sky130_fd_sc_hd__a21o_1 _379_ (.A1(_060_),
    .A2(_061_),
    .B1(_038_),
    .X(_063_));
 sky130_fd_sc_hd__nand2b_1 _380_ (.A_N(_062_),
    .B(_063_),
    .Y(_064_));
 sky130_fd_sc_hd__xnor2_1 _381_ (.A(_040_),
    .B(_064_),
    .Y(\Adder.cla_16_bit.Sum[4] ));
 sky130_fd_sc_hd__or2_1 _382_ (.A(_043_),
    .B(_044_),
    .X(_065_));
 sky130_fd_sc_hd__or3b_2 _383_ (.A(\B_ff[3] ),
    .B(\B_ff[4] ),
    .C_N(\B_ff[5] ),
    .X(_066_));
 sky130_fd_sc_hd__or3_1 _384_ (.A(_283_),
    .B(\B_ff[5] ),
    .C(_042_),
    .X(_067_));
 sky130_fd_sc_hd__nor2_2 _385_ (.A(_041_),
    .B(_046_),
    .Y(_068_));
 sky130_fd_sc_hd__nand2_1 _386_ (.A(_042_),
    .B(_045_),
    .Y(_069_));
 sky130_fd_sc_hd__o221a_1 _387_ (.A1(\A_ff[1] ),
    .A2(_065_),
    .B1(_066_),
    .B2(\A_ff[0] ),
    .C1(_067_),
    .X(_070_));
 sky130_fd_sc_hd__a21bo_1 _388_ (.A1(\A_ff[1] ),
    .A2(_068_),
    .B1_N(_070_),
    .X(_071_));
 sky130_fd_sc_hd__nor2_1 _389_ (.A(\A_ff[4] ),
    .B(_292_),
    .Y(_072_));
 sky130_fd_sc_hd__mux2_1 _390_ (.A0(_290_),
    .A1(_293_),
    .S(\A_ff[5] ),
    .X(_073_));
 sky130_fd_sc_hd__nor2_1 _391_ (.A(_072_),
    .B(_073_),
    .Y(_074_));
 sky130_fd_sc_hd__o21ai_1 _392_ (.A1(\A_ff[2] ),
    .A2(_298_),
    .B1(_311_),
    .Y(_075_));
 sky130_fd_sc_hd__o22a_1 _393_ (.A1(\A_ff[3] ),
    .A2(_299_),
    .B1(_306_),
    .B2(\A_ff[2] ),
    .X(_076_));
 sky130_fd_sc_hd__o2bb2a_1 _394_ (.A1_N(_075_),
    .A2_N(_076_),
    .B1(\A_ff[3] ),
    .B2(_032_),
    .X(_077_));
 sky130_fd_sc_hd__and2b_1 _395_ (.A_N(_074_),
    .B(_077_),
    .X(_078_));
 sky130_fd_sc_hd__or3_1 _396_ (.A(_072_),
    .B(_073_),
    .C(_077_),
    .X(_079_));
 sky130_fd_sc_hd__xnor2_1 _397_ (.A(_074_),
    .B(_077_),
    .Y(_080_));
 sky130_fd_sc_hd__o21ai_2 _398_ (.A1(_071_),
    .A2(_078_),
    .B1(_079_),
    .Y(_081_));
 sky130_fd_sc_hd__xnor2_1 _399_ (.A(_071_),
    .B(_080_),
    .Y(_082_));
 sky130_fd_sc_hd__a21bo_1 _400_ (.A1(_049_),
    .A2(_057_),
    .B1_N(_056_),
    .X(_083_));
 sky130_fd_sc_hd__nand2b_1 _401_ (.A_N(_082_),
    .B(_083_),
    .Y(_084_));
 sky130_fd_sc_hd__xnor2_1 _402_ (.A(_082_),
    .B(_083_),
    .Y(_085_));
 sky130_fd_sc_hd__and2b_1 _403_ (.A_N(_060_),
    .B(_085_),
    .X(_086_));
 sky130_fd_sc_hd__xnor2_1 _404_ (.A(_060_),
    .B(_085_),
    .Y(_087_));
 sky130_fd_sc_hd__a21o_1 _405_ (.A1(_040_),
    .A2(_063_),
    .B1(_062_),
    .X(_088_));
 sky130_fd_sc_hd__xor2_1 _406_ (.A(_087_),
    .B(_088_),
    .X(\Adder.cla_16_bit.Sum[5] ));
 sky130_fd_sc_hd__and2_1 _407_ (.A(\B_ff[5] ),
    .B(\B_ff[6] ),
    .X(_089_));
 sky130_fd_sc_hd__nand2_1 _408_ (.A(\B_ff[5] ),
    .B(\B_ff[6] ),
    .Y(_090_));
 sky130_fd_sc_hd__nor2_1 _409_ (.A(\B_ff[5] ),
    .B(\B_ff[6] ),
    .Y(_091_));
 sky130_fd_sc_hd__and3b_1 _410_ (.A_N(_091_),
    .B(\A_ff[0] ),
    .C(_090_),
    .X(_092_));
 sky130_fd_sc_hd__o21ai_1 _411_ (.A1(\A_ff[1] ),
    .A2(_042_),
    .B1(_045_),
    .Y(_093_));
 sky130_fd_sc_hd__o221a_1 _412_ (.A1(\A_ff[2] ),
    .A2(_065_),
    .B1(_066_),
    .B2(\A_ff[1] ),
    .C1(_093_),
    .X(_094_));
 sky130_fd_sc_hd__a21oi_1 _413_ (.A1(_284_),
    .A2(_068_),
    .B1(_094_),
    .Y(_095_));
 sky130_fd_sc_hd__mux2_1 _414_ (.A0(_291_),
    .A1(_294_),
    .S(\A_ff[6] ),
    .X(_096_));
 sky130_fd_sc_hd__o21ai_1 _415_ (.A1(\A_ff[5] ),
    .A2(_292_),
    .B1(_096_),
    .Y(_097_));
 sky130_fd_sc_hd__o21ai_1 _416_ (.A1(\A_ff[3] ),
    .A2(_298_),
    .B1(_311_),
    .Y(_098_));
 sky130_fd_sc_hd__o22a_1 _417_ (.A1(\A_ff[4] ),
    .A2(_299_),
    .B1(_306_),
    .B2(\A_ff[3] ),
    .X(_099_));
 sky130_fd_sc_hd__o2bb2a_1 _418_ (.A1_N(_098_),
    .A2_N(_099_),
    .B1(\A_ff[4] ),
    .B2(_032_),
    .X(_100_));
 sky130_fd_sc_hd__and2_1 _419_ (.A(_097_),
    .B(_100_),
    .X(_101_));
 sky130_fd_sc_hd__or2_1 _420_ (.A(_097_),
    .B(_100_),
    .X(_102_));
 sky130_fd_sc_hd__xor2_1 _421_ (.A(_097_),
    .B(_100_),
    .X(_103_));
 sky130_fd_sc_hd__xnor2_1 _422_ (.A(_095_),
    .B(_103_),
    .Y(_104_));
 sky130_fd_sc_hd__and2b_1 _423_ (.A_N(_092_),
    .B(_104_),
    .X(_105_));
 sky130_fd_sc_hd__nand2b_1 _424_ (.A_N(_104_),
    .B(_092_),
    .Y(_106_));
 sky130_fd_sc_hd__xor2_1 _425_ (.A(_092_),
    .B(_104_),
    .X(_107_));
 sky130_fd_sc_hd__a21o_1 _426_ (.A1(_081_),
    .A2(_106_),
    .B1(_105_),
    .X(_108_));
 sky130_fd_sc_hd__xnor2_2 _427_ (.A(_081_),
    .B(_107_),
    .Y(_109_));
 sky130_fd_sc_hd__nor2_1 _428_ (.A(_084_),
    .B(_109_),
    .Y(_110_));
 sky130_fd_sc_hd__xor2_1 _429_ (.A(_084_),
    .B(_109_),
    .X(_111_));
 sky130_fd_sc_hd__a21o_1 _430_ (.A1(_087_),
    .A2(_088_),
    .B1(_086_),
    .X(_112_));
 sky130_fd_sc_hd__xor2_1 _431_ (.A(_111_),
    .B(_112_),
    .X(\Adder.cla_16_bit.Sum[6] ));
 sky130_fd_sc_hd__a21o_1 _432_ (.A1(_111_),
    .A2(_112_),
    .B1(_110_),
    .X(_113_));
 sky130_fd_sc_hd__nand2_2 _433_ (.A(\B_ff[7] ),
    .B(_091_),
    .Y(_114_));
 sky130_fd_sc_hd__nor2_1 _434_ (.A(\B_ff[7] ),
    .B(_090_),
    .Y(_115_));
 sky130_fd_sc_hd__nor2_1 _435_ (.A(_283_),
    .B(_115_),
    .Y(_116_));
 sky130_fd_sc_hd__a21oi_1 _436_ (.A1(_283_),
    .A2(_114_),
    .B1(_116_),
    .Y(_117_));
 sky130_fd_sc_hd__nor2_1 _437_ (.A(\B_ff[7] ),
    .B(_091_),
    .Y(_118_));
 sky130_fd_sc_hd__or2_1 _438_ (.A(\B_ff[7] ),
    .B(_091_),
    .X(_119_));
 sky130_fd_sc_hd__nor2_1 _439_ (.A(_089_),
    .B(_119_),
    .Y(_120_));
 sky130_fd_sc_hd__nand2_1 _440_ (.A(_090_),
    .B(_118_),
    .Y(_121_));
 sky130_fd_sc_hd__nand2_1 _441_ (.A(\B_ff[7] ),
    .B(_090_),
    .Y(_122_));
 sky130_fd_sc_hd__or2_2 _442_ (.A(_091_),
    .B(_122_),
    .X(_123_));
 sky130_fd_sc_hd__nor2_1 _443_ (.A(\A_ff[1] ),
    .B(_123_),
    .Y(_124_));
 sky130_fd_sc_hd__a211o_1 _444_ (.A1(\A_ff[1] ),
    .A2(_120_),
    .B1(_124_),
    .C1(_117_),
    .X(_125_));
 sky130_fd_sc_hd__o21a_1 _445_ (.A1(_095_),
    .A2(_101_),
    .B1(_102_),
    .X(_126_));
 sky130_fd_sc_hd__nor2_1 _446_ (.A(\A_ff[6] ),
    .B(_292_),
    .Y(_127_));
 sky130_fd_sc_hd__mux2_1 _447_ (.A0(_290_),
    .A1(_293_),
    .S(\A_ff[7] ),
    .X(_128_));
 sky130_fd_sc_hd__nor2_1 _448_ (.A(_127_),
    .B(_128_),
    .Y(_129_));
 sky130_fd_sc_hd__mux2_1 _449_ (.A0(_305_),
    .A1(_311_),
    .S(\A_ff[4] ),
    .X(_130_));
 sky130_fd_sc_hd__a21oi_1 _450_ (.A1(\B_ff[3] ),
    .A2(\A_ff[5] ),
    .B1(_299_),
    .Y(_131_));
 sky130_fd_sc_hd__o22a_1 _451_ (.A1(\A_ff[5] ),
    .A2(_032_),
    .B1(_130_),
    .B2(_131_),
    .X(_132_));
 sky130_fd_sc_hd__or3_1 _452_ (.A(_127_),
    .B(_128_),
    .C(_132_),
    .X(_133_));
 sky130_fd_sc_hd__and2b_1 _453_ (.A_N(_129_),
    .B(_132_),
    .X(_134_));
 sky130_fd_sc_hd__xnor2_1 _454_ (.A(_129_),
    .B(_132_),
    .Y(_135_));
 sky130_fd_sc_hd__nor2_1 _455_ (.A(\A_ff[3] ),
    .B(_065_),
    .Y(_136_));
 sky130_fd_sc_hd__nor2_1 _456_ (.A(\A_ff[2] ),
    .B(_066_),
    .Y(_137_));
 sky130_fd_sc_hd__a21oi_1 _457_ (.A1(_284_),
    .A2(_041_),
    .B1(_046_),
    .Y(_138_));
 sky130_fd_sc_hd__o32a_1 _458_ (.A1(_136_),
    .A2(_137_),
    .A3(_138_),
    .B1(_069_),
    .B2(\A_ff[3] ),
    .X(_139_));
 sky130_fd_sc_hd__xnor2_1 _459_ (.A(_135_),
    .B(_139_),
    .Y(_140_));
 sky130_fd_sc_hd__nand2b_1 _460_ (.A_N(_126_),
    .B(_140_),
    .Y(_141_));
 sky130_fd_sc_hd__and2b_1 _461_ (.A_N(_140_),
    .B(_126_),
    .X(_142_));
 sky130_fd_sc_hd__xnor2_1 _462_ (.A(_126_),
    .B(_140_),
    .Y(_143_));
 sky130_fd_sc_hd__o21ai_1 _463_ (.A1(\A_ff[0] ),
    .A2(_123_),
    .B1(_114_),
    .Y(_144_));
 sky130_fd_sc_hd__xnor2_1 _464_ (.A(_143_),
    .B(_144_),
    .Y(_145_));
 sky130_fd_sc_hd__nand2_1 _465_ (.A(_108_),
    .B(_145_),
    .Y(_146_));
 sky130_fd_sc_hd__xnor2_1 _466_ (.A(_108_),
    .B(_145_),
    .Y(_147_));
 sky130_fd_sc_hd__o21bai_1 _467_ (.A1(_108_),
    .A2(_145_),
    .B1_N(_125_),
    .Y(_148_));
 sky130_fd_sc_hd__xnor2_2 _468_ (.A(_125_),
    .B(_147_),
    .Y(_149_));
 sky130_fd_sc_hd__xor2_1 _469_ (.A(_113_),
    .B(_149_),
    .X(\Adder.cla_16_bit.Sum[7] ));
 sky130_fd_sc_hd__nand2_1 _470_ (.A(\A_ff[1] ),
    .B(_115_),
    .Y(_150_));
 sky130_fd_sc_hd__o221a_1 _471_ (.A1(\A_ff[1] ),
    .A2(_114_),
    .B1(_123_),
    .B2(\A_ff[2] ),
    .C1(_150_),
    .X(_151_));
 sky130_fd_sc_hd__o21ai_1 _472_ (.A1(_284_),
    .A2(_121_),
    .B1(_151_),
    .Y(_152_));
 sky130_fd_sc_hd__o21ai_1 _473_ (.A1(\A_ff[3] ),
    .A2(_042_),
    .B1(_045_),
    .Y(_153_));
 sky130_fd_sc_hd__o221a_1 _474_ (.A1(\A_ff[4] ),
    .A2(_065_),
    .B1(_066_),
    .B2(\A_ff[3] ),
    .C1(_153_),
    .X(_154_));
 sky130_fd_sc_hd__a21oi_2 _475_ (.A1(_285_),
    .A2(_068_),
    .B1(_154_),
    .Y(_155_));
 sky130_fd_sc_hd__mux2_2 _476_ (.A0(\B_ff[1] ),
    .A1(_293_),
    .S(\A_ff[7] ),
    .X(_156_));
 sky130_fd_sc_hd__mux2_1 _477_ (.A0(_305_),
    .A1(_311_),
    .S(\A_ff[5] ),
    .X(_157_));
 sky130_fd_sc_hd__a21oi_1 _478_ (.A1(\B_ff[3] ),
    .A2(\A_ff[6] ),
    .B1(_299_),
    .Y(_158_));
 sky130_fd_sc_hd__o22a_1 _479_ (.A1(\A_ff[6] ),
    .A2(_032_),
    .B1(_157_),
    .B2(_158_),
    .X(_159_));
 sky130_fd_sc_hd__and2_1 _480_ (.A(_156_),
    .B(_159_),
    .X(_160_));
 sky130_fd_sc_hd__or2_1 _481_ (.A(_156_),
    .B(_159_),
    .X(_161_));
 sky130_fd_sc_hd__xnor2_1 _482_ (.A(_156_),
    .B(_159_),
    .Y(_162_));
 sky130_fd_sc_hd__xnor2_1 _483_ (.A(_155_),
    .B(_162_),
    .Y(_163_));
 sky130_fd_sc_hd__a21o_1 _484_ (.A1(_133_),
    .A2(_139_),
    .B1(_134_),
    .X(_164_));
 sky130_fd_sc_hd__xor2_1 _485_ (.A(_163_),
    .B(_164_),
    .X(_165_));
 sky130_fd_sc_hd__o21a_1 _486_ (.A1(_163_),
    .A2(_164_),
    .B1(_152_),
    .X(_166_));
 sky130_fd_sc_hd__a21oi_1 _487_ (.A1(_163_),
    .A2(_164_),
    .B1(_166_),
    .Y(_167_));
 sky130_fd_sc_hd__xnor2_1 _488_ (.A(_152_),
    .B(_165_),
    .Y(_168_));
 sky130_fd_sc_hd__a21oi_1 _489_ (.A1(_141_),
    .A2(_144_),
    .B1(_142_),
    .Y(_169_));
 sky130_fd_sc_hd__nor2_1 _490_ (.A(_168_),
    .B(_169_),
    .Y(_170_));
 sky130_fd_sc_hd__xor2_1 _491_ (.A(_168_),
    .B(_169_),
    .X(_171_));
 sky130_fd_sc_hd__a21o_1 _492_ (.A1(_146_),
    .A2(_148_),
    .B1(_171_),
    .X(_172_));
 sky130_fd_sc_hd__and3_1 _493_ (.A(_146_),
    .B(_148_),
    .C(_171_),
    .X(_173_));
 sky130_fd_sc_hd__nand3_1 _494_ (.A(_146_),
    .B(_148_),
    .C(_171_),
    .Y(_174_));
 sky130_fd_sc_hd__and4_1 _495_ (.A(_113_),
    .B(_149_),
    .C(_172_),
    .D(_174_),
    .X(_175_));
 sky130_fd_sc_hd__a22o_1 _496_ (.A1(_113_),
    .A2(_149_),
    .B1(_172_),
    .B2(_174_),
    .X(_176_));
 sky130_fd_sc_hd__and2b_1 _497_ (.A_N(_175_),
    .B(_176_),
    .X(\Adder.cla_16_bit.Sum[8] ));
 sky130_fd_sc_hd__nand2_1 _498_ (.A(\A_ff[2] ),
    .B(_115_),
    .Y(_177_));
 sky130_fd_sc_hd__o221a_1 _499_ (.A1(\A_ff[2] ),
    .A2(_114_),
    .B1(_123_),
    .B2(\A_ff[3] ),
    .C1(_177_),
    .X(_178_));
 sky130_fd_sc_hd__a21bo_1 _500_ (.A1(\A_ff[3] ),
    .A2(_120_),
    .B1_N(_178_),
    .X(_179_));
 sky130_fd_sc_hd__o21ai_2 _501_ (.A1(_155_),
    .A2(_160_),
    .B1(_161_),
    .Y(_180_));
 sky130_fd_sc_hd__mux2_1 _502_ (.A0(_305_),
    .A1(_311_),
    .S(\A_ff[6] ),
    .X(_181_));
 sky130_fd_sc_hd__a21oi_1 _503_ (.A1(\B_ff[3] ),
    .A2(\A_ff[7] ),
    .B1(_299_),
    .Y(_182_));
 sky130_fd_sc_hd__o22a_1 _504_ (.A1(\A_ff[7] ),
    .A2(_032_),
    .B1(_181_),
    .B2(_182_),
    .X(_183_));
 sky130_fd_sc_hd__xor2_1 _505_ (.A(_156_),
    .B(_183_),
    .X(_184_));
 sky130_fd_sc_hd__mux2_1 _506_ (.A0(_046_),
    .A1(_066_),
    .S(_285_),
    .X(_185_));
 sky130_fd_sc_hd__a211o_1 _507_ (.A1(\B_ff[5] ),
    .A2(\A_ff[5] ),
    .B1(_041_),
    .C1(_044_),
    .X(_186_));
 sky130_fd_sc_hd__o2bb2a_1 _508_ (.A1_N(_186_),
    .A2_N(_185_),
    .B1(_069_),
    .B2(\A_ff[5] ),
    .X(_187_));
 sky130_fd_sc_hd__xnor2_1 _509_ (.A(_184_),
    .B(_187_),
    .Y(_188_));
 sky130_fd_sc_hd__xor2_1 _510_ (.A(_180_),
    .B(_188_),
    .X(_189_));
 sky130_fd_sc_hd__o21ba_1 _511_ (.A1(_180_),
    .A2(_188_),
    .B1_N(_179_),
    .X(_190_));
 sky130_fd_sc_hd__a21o_1 _512_ (.A1(_180_),
    .A2(_188_),
    .B1(_190_),
    .X(_191_));
 sky130_fd_sc_hd__xnor2_1 _513_ (.A(_179_),
    .B(_189_),
    .Y(_192_));
 sky130_fd_sc_hd__nor2_1 _514_ (.A(_167_),
    .B(_192_),
    .Y(_193_));
 sky130_fd_sc_hd__xor2_1 _515_ (.A(_167_),
    .B(_192_),
    .X(_194_));
 sky130_fd_sc_hd__nand2_1 _516_ (.A(_170_),
    .B(_194_),
    .Y(_195_));
 sky130_fd_sc_hd__xnor2_1 _517_ (.A(_170_),
    .B(_194_),
    .Y(_196_));
 sky130_fd_sc_hd__inv_2 _518_ (.A(_196_),
    .Y(_197_));
 sky130_fd_sc_hd__a31o_1 _519_ (.A1(_113_),
    .A2(_149_),
    .A3(_172_),
    .B1(_173_),
    .X(_198_));
 sky130_fd_sc_hd__nand2_1 _520_ (.A(_197_),
    .B(_198_),
    .Y(_199_));
 sky130_fd_sc_hd__xnor2_1 _521_ (.A(_196_),
    .B(_198_),
    .Y(\Adder.cla_16_bit.Sum[9] ));
 sky130_fd_sc_hd__mux2_1 _522_ (.A0(_303_),
    .A1(_311_),
    .S(\A_ff[7] ),
    .X(_200_));
 sky130_fd_sc_hd__and2_1 _523_ (.A(_156_),
    .B(_200_),
    .X(_201_));
 sky130_fd_sc_hd__or3_1 _524_ (.A(\A_ff[6] ),
    .B(_043_),
    .C(_044_),
    .X(_202_));
 sky130_fd_sc_hd__or2_1 _525_ (.A(\A_ff[5] ),
    .B(_066_),
    .X(_203_));
 sky130_fd_sc_hd__o21ai_1 _526_ (.A1(\A_ff[5] ),
    .A2(_042_),
    .B1(_045_),
    .Y(_204_));
 sky130_fd_sc_hd__a32o_1 _527_ (.A1(_202_),
    .A2(_203_),
    .A3(_204_),
    .B1(_068_),
    .B2(_286_),
    .X(_205_));
 sky130_fd_sc_hd__nor2_1 _528_ (.A(_156_),
    .B(_200_),
    .Y(_206_));
 sky130_fd_sc_hd__nor2_1 _529_ (.A(_205_),
    .B(_206_),
    .Y(_207_));
 sky130_fd_sc_hd__xnor2_1 _530_ (.A(_156_),
    .B(_200_),
    .Y(_208_));
 sky130_fd_sc_hd__xnor2_1 _531_ (.A(_205_),
    .B(_208_),
    .Y(_209_));
 sky130_fd_sc_hd__o21a_1 _532_ (.A1(_156_),
    .A2(_183_),
    .B1(_187_),
    .X(_210_));
 sky130_fd_sc_hd__a21oi_1 _533_ (.A1(_156_),
    .A2(_183_),
    .B1(_210_),
    .Y(_211_));
 sky130_fd_sc_hd__xnor2_1 _534_ (.A(_209_),
    .B(_211_),
    .Y(_212_));
 sky130_fd_sc_hd__nand2_1 _535_ (.A(\A_ff[3] ),
    .B(_115_),
    .Y(_213_));
 sky130_fd_sc_hd__o221a_1 _536_ (.A1(\A_ff[3] ),
    .A2(_114_),
    .B1(_123_),
    .B2(\A_ff[4] ),
    .C1(_213_),
    .X(_214_));
 sky130_fd_sc_hd__mux2_1 _537_ (.A0(_285_),
    .A1(_214_),
    .S(_121_),
    .X(_215_));
 sky130_fd_sc_hd__xor2_1 _538_ (.A(_212_),
    .B(_215_),
    .X(_216_));
 sky130_fd_sc_hd__and2b_1 _539_ (.A_N(_191_),
    .B(_216_),
    .X(_217_));
 sky130_fd_sc_hd__xnor2_1 _540_ (.A(_191_),
    .B(_216_),
    .Y(_218_));
 sky130_fd_sc_hd__nor2_1 _541_ (.A(_193_),
    .B(_218_),
    .Y(_219_));
 sky130_fd_sc_hd__nand2_1 _542_ (.A(_193_),
    .B(_218_),
    .Y(_220_));
 sky130_fd_sc_hd__nand2b_1 _543_ (.A_N(_219_),
    .B(_220_),
    .Y(_221_));
 sky130_fd_sc_hd__a21o_1 _544_ (.A1(_195_),
    .A2(_199_),
    .B1(_221_),
    .X(_222_));
 sky130_fd_sc_hd__and2_1 _545_ (.A(_199_),
    .B(_221_),
    .X(_223_));
 sky130_fd_sc_hd__a21boi_1 _546_ (.A1(_195_),
    .A2(_223_),
    .B1_N(_222_),
    .Y(\Adder.cla_16_bit.Sum[10] ));
 sky130_fd_sc_hd__nand2_1 _547_ (.A(_220_),
    .B(_222_),
    .Y(_224_));
 sky130_fd_sc_hd__o21a_1 _548_ (.A1(_209_),
    .A2(_211_),
    .B1(_215_),
    .X(_225_));
 sky130_fd_sc_hd__a21oi_1 _549_ (.A1(_209_),
    .A2(_211_),
    .B1(_225_),
    .Y(_226_));
 sky130_fd_sc_hd__or3_1 _550_ (.A(\A_ff[7] ),
    .B(_043_),
    .C(_044_),
    .X(_227_));
 sky130_fd_sc_hd__or2_1 _551_ (.A(\A_ff[6] ),
    .B(_066_),
    .X(_228_));
 sky130_fd_sc_hd__a21o_1 _552_ (.A1(_286_),
    .A2(_041_),
    .B1(_046_),
    .X(_229_));
 sky130_fd_sc_hd__a32oi_4 _553_ (.A1(_227_),
    .A2(_228_),
    .A3(_229_),
    .B1(_068_),
    .B2(_287_),
    .Y(_230_));
 sky130_fd_sc_hd__nor2_1 _554_ (.A(_206_),
    .B(_230_),
    .Y(_231_));
 sky130_fd_sc_hd__xnor2_1 _555_ (.A(_208_),
    .B(_230_),
    .Y(_232_));
 sky130_fd_sc_hd__o21ai_1 _556_ (.A1(_201_),
    .A2(_207_),
    .B1(_232_),
    .Y(_233_));
 sky130_fd_sc_hd__or3_1 _557_ (.A(_201_),
    .B(_207_),
    .C(_232_),
    .X(_234_));
 sky130_fd_sc_hd__nand2_1 _558_ (.A(_233_),
    .B(_234_),
    .Y(_235_));
 sky130_fd_sc_hd__a21o_1 _559_ (.A1(_285_),
    .A2(_089_),
    .B1(_119_),
    .X(_236_));
 sky130_fd_sc_hd__o221a_1 _560_ (.A1(\A_ff[4] ),
    .A2(_114_),
    .B1(_123_),
    .B2(\A_ff[5] ),
    .C1(_236_),
    .X(_237_));
 sky130_fd_sc_hd__o21ba_1 _561_ (.A1(\A_ff[5] ),
    .A2(_121_),
    .B1_N(_237_),
    .X(_238_));
 sky130_fd_sc_hd__xor2_1 _562_ (.A(_235_),
    .B(_238_),
    .X(_239_));
 sky130_fd_sc_hd__nand2b_1 _563_ (.A_N(_239_),
    .B(_226_),
    .Y(_240_));
 sky130_fd_sc_hd__xnor2_1 _564_ (.A(_226_),
    .B(_239_),
    .Y(_241_));
 sky130_fd_sc_hd__nor2_1 _565_ (.A(_217_),
    .B(_241_),
    .Y(_242_));
 sky130_fd_sc_hd__nand2_1 _566_ (.A(_217_),
    .B(_241_),
    .Y(_243_));
 sky130_fd_sc_hd__nand2b_1 _567_ (.A_N(_242_),
    .B(_243_),
    .Y(_244_));
 sky130_fd_sc_hd__xnor2_1 _568_ (.A(_224_),
    .B(_244_),
    .Y(\Adder.cla_16_bit.Sum[11] ));
 sky130_fd_sc_hd__o21ai_1 _569_ (.A1(\A_ff[5] ),
    .A2(_090_),
    .B1(_118_),
    .Y(_245_));
 sky130_fd_sc_hd__o221a_1 _570_ (.A1(\A_ff[5] ),
    .A2(_114_),
    .B1(_123_),
    .B2(\A_ff[6] ),
    .C1(_245_),
    .X(_246_));
 sky130_fd_sc_hd__a21oi_1 _571_ (.A1(_286_),
    .A2(_120_),
    .B1(_246_),
    .Y(_247_));
 sky130_fd_sc_hd__mux2_1 _572_ (.A0(_043_),
    .A1(_046_),
    .S(\A_ff[7] ),
    .X(_248_));
 sky130_fd_sc_hd__nand2_1 _573_ (.A(_247_),
    .B(_248_),
    .Y(_249_));
 sky130_fd_sc_hd__xor2_1 _574_ (.A(_247_),
    .B(_248_),
    .X(_250_));
 sky130_fd_sc_hd__nor2_1 _575_ (.A(_201_),
    .B(_231_),
    .Y(_251_));
 sky130_fd_sc_hd__xor2_1 _576_ (.A(_250_),
    .B(_251_),
    .X(_252_));
 sky130_fd_sc_hd__a21bo_1 _577_ (.A1(_234_),
    .A2(_238_),
    .B1_N(_233_),
    .X(_253_));
 sky130_fd_sc_hd__and2_1 _578_ (.A(_252_),
    .B(_253_),
    .X(_254_));
 sky130_fd_sc_hd__nor2_1 _579_ (.A(_252_),
    .B(_253_),
    .Y(_255_));
 sky130_fd_sc_hd__or2_1 _580_ (.A(_254_),
    .B(_255_),
    .X(_256_));
 sky130_fd_sc_hd__nor2_1 _581_ (.A(_240_),
    .B(_256_),
    .Y(_257_));
 sky130_fd_sc_hd__and2_1 _582_ (.A(_240_),
    .B(_256_),
    .X(_258_));
 sky130_fd_sc_hd__nor2_1 _583_ (.A(_257_),
    .B(_258_),
    .Y(_259_));
 sky130_fd_sc_hd__o211a_1 _584_ (.A1(_220_),
    .A2(_242_),
    .B1(_243_),
    .C1(_195_),
    .X(_260_));
 sky130_fd_sc_hd__a21bo_1 _585_ (.A1(_197_),
    .A2(_198_),
    .B1_N(_260_),
    .X(_261_));
 sky130_fd_sc_hd__o21ai_1 _586_ (.A1(_219_),
    .A2(_242_),
    .B1(_243_),
    .Y(_262_));
 sky130_fd_sc_hd__and3_1 _587_ (.A(_259_),
    .B(_261_),
    .C(_262_),
    .X(_263_));
 sky130_fd_sc_hd__a21oi_1 _588_ (.A1(_261_),
    .A2(_262_),
    .B1(_259_),
    .Y(_264_));
 sky130_fd_sc_hd__nor2_1 _589_ (.A(_263_),
    .B(_264_),
    .Y(\Adder.cla_16_bit.Sum[12] ));
 sky130_fd_sc_hd__nand2_1 _590_ (.A(\A_ff[6] ),
    .B(_115_),
    .Y(_265_));
 sky130_fd_sc_hd__o221a_1 _591_ (.A1(\A_ff[6] ),
    .A2(_114_),
    .B1(_123_),
    .B2(\A_ff[7] ),
    .C1(_121_),
    .X(_266_));
 sky130_fd_sc_hd__a22o_1 _592_ (.A1(_287_),
    .A2(_120_),
    .B1(_265_),
    .B2(_266_),
    .X(_267_));
 sky130_fd_sc_hd__and3_1 _593_ (.A(_250_),
    .B(_251_),
    .C(_267_),
    .X(_268_));
 sky130_fd_sc_hd__nand2_1 _594_ (.A(_249_),
    .B(_267_),
    .Y(_269_));
 sky130_fd_sc_hd__o2bb2a_1 _595_ (.A1_N(_250_),
    .A2_N(_251_),
    .B1(_267_),
    .B2(_249_),
    .X(_270_));
 sky130_fd_sc_hd__a21oi_1 _596_ (.A1(_269_),
    .A2(_270_),
    .B1(_268_),
    .Y(_271_));
 sky130_fd_sc_hd__and2_1 _597_ (.A(_254_),
    .B(_271_),
    .X(_272_));
 sky130_fd_sc_hd__or2_1 _598_ (.A(_254_),
    .B(_271_),
    .X(_273_));
 sky130_fd_sc_hd__nand2b_1 _599_ (.A_N(_272_),
    .B(_273_),
    .Y(_274_));
 sky130_fd_sc_hd__a31o_1 _600_ (.A1(_259_),
    .A2(_261_),
    .A3(_262_),
    .B1(_257_),
    .X(_275_));
 sky130_fd_sc_hd__xnor2_1 _601_ (.A(_274_),
    .B(_275_),
    .Y(\Adder.cla_16_bit.Sum[13] ));
 sky130_fd_sc_hd__mux2_1 _602_ (.A0(_119_),
    .A1(_122_),
    .S(_287_),
    .X(_276_));
 sky130_fd_sc_hd__or2_1 _603_ (.A(_269_),
    .B(_276_),
    .X(_277_));
 sky130_fd_sc_hd__nand2_1 _604_ (.A(_269_),
    .B(_276_),
    .Y(_278_));
 sky130_fd_sc_hd__and2_1 _605_ (.A(_277_),
    .B(_278_),
    .X(_279_));
 sky130_fd_sc_hd__nand2_1 _606_ (.A(_268_),
    .B(_279_),
    .Y(_280_));
 sky130_fd_sc_hd__xnor2_1 _607_ (.A(_268_),
    .B(_279_),
    .Y(_281_));
 sky130_fd_sc_hd__a21oi_1 _608_ (.A1(_273_),
    .A2(_275_),
    .B1(_272_),
    .Y(_282_));
 sky130_fd_sc_hd__xor2_1 _609_ (.A(_281_),
    .B(_282_),
    .X(\Adder.cla_16_bit.Sum[14] ));
 sky130_fd_sc_hd__o211a_1 _610_ (.A1(_281_),
    .A2(_282_),
    .B1(_278_),
    .C1(_280_),
    .X(\Adder.cla_16_bit.Sum[15] ));
 sky130_fd_sc_hd__inv_2 _611_ (.A(net17),
    .Y(_001_));
 sky130_fd_sc_hd__inv_2 _612_ (.A(net17),
    .Y(_002_));
 sky130_fd_sc_hd__inv_2 _613_ (.A(net17),
    .Y(_003_));
 sky130_fd_sc_hd__inv_2 _614_ (.A(net17),
    .Y(_004_));
 sky130_fd_sc_hd__inv_2 _615_ (.A(net17),
    .Y(_005_));
 sky130_fd_sc_hd__inv_2 _616_ (.A(net17),
    .Y(_006_));
 sky130_fd_sc_hd__inv_2 _617_ (.A(net17),
    .Y(_007_));
 sky130_fd_sc_hd__inv_2 _618_ (.A(net17),
    .Y(_008_));
 sky130_fd_sc_hd__inv_2 _619_ (.A(net17),
    .Y(_009_));
 sky130_fd_sc_hd__inv_2 _620_ (.A(net17),
    .Y(_010_));
 sky130_fd_sc_hd__inv_2 _621_ (.A(net17),
    .Y(_011_));
 sky130_fd_sc_hd__inv_2 _622_ (.A(net17),
    .Y(_012_));
 sky130_fd_sc_hd__inv_2 _623_ (.A(net17),
    .Y(_013_));
 sky130_fd_sc_hd__inv_2 _624_ (.A(net17),
    .Y(_014_));
 sky130_fd_sc_hd__inv_2 _625_ (.A(net17),
    .Y(_015_));
 sky130_fd_sc_hd__inv_2 _626_ (.A(net17),
    .Y(_016_));
 sky130_fd_sc_hd__inv_2 _627_ (.A(net17),
    .Y(_017_));
 sky130_fd_sc_hd__inv_2 _628_ (.A(net17),
    .Y(_018_));
 sky130_fd_sc_hd__inv_2 _629_ (.A(net17),
    .Y(_019_));
 sky130_fd_sc_hd__inv_2 _630_ (.A(net17),
    .Y(_020_));
 sky130_fd_sc_hd__inv_2 _631_ (.A(net17),
    .Y(_021_));
 sky130_fd_sc_hd__inv_2 _632_ (.A(net17),
    .Y(_022_));
 sky130_fd_sc_hd__inv_2 _633_ (.A(net17),
    .Y(_023_));
 sky130_fd_sc_hd__inv_2 _634_ (.A(net17),
    .Y(_024_));
 sky130_fd_sc_hd__inv_2 _635_ (.A(net17),
    .Y(_025_));
 sky130_fd_sc_hd__inv_2 _636_ (.A(net17),
    .Y(_026_));
 sky130_fd_sc_hd__inv_2 _637_ (.A(net17),
    .Y(_027_));
 sky130_fd_sc_hd__inv_2 _638_ (.A(net17),
    .Y(_028_));
 sky130_fd_sc_hd__inv_2 _639_ (.A(net17),
    .Y(_029_));
 sky130_fd_sc_hd__inv_2 _640_ (.A(net17),
    .Y(_030_));
 sky130_fd_sc_hd__inv_2 _641_ (.A(net17),
    .Y(_031_));
 sky130_fd_sc_hd__dfrtp_1 _642_ (.CLK(clknet_2_0__leaf_clk),
    .D(\Adder.cla_16_bit.Sum[0] ),
    .RESET_B(_000_),
    .Q(net18));
 sky130_fd_sc_hd__dfrtp_1 _643_ (.CLK(clknet_2_0__leaf_clk),
    .D(\Adder.cla_16_bit.Sum[1] ),
    .RESET_B(_001_),
    .Q(net25));
 sky130_fd_sc_hd__dfrtp_1 _644_ (.CLK(clknet_2_0__leaf_clk),
    .D(\Adder.cla_16_bit.Sum[2] ),
    .RESET_B(_002_),
    .Q(net26));
 sky130_fd_sc_hd__dfrtp_1 _645_ (.CLK(clknet_2_0__leaf_clk),
    .D(\Adder.cla_16_bit.Sum[3] ),
    .RESET_B(_003_),
    .Q(net27));
 sky130_fd_sc_hd__dfrtp_1 _646_ (.CLK(clknet_2_0__leaf_clk),
    .D(\Adder.cla_16_bit.Sum[4] ),
    .RESET_B(_004_),
    .Q(net28));
 sky130_fd_sc_hd__dfrtp_1 _647_ (.CLK(clknet_2_0__leaf_clk),
    .D(\Adder.cla_16_bit.Sum[5] ),
    .RESET_B(_005_),
    .Q(net29));
 sky130_fd_sc_hd__dfrtp_1 _648_ (.CLK(clknet_2_0__leaf_clk),
    .D(\Adder.cla_16_bit.Sum[6] ),
    .RESET_B(_006_),
    .Q(net30));
 sky130_fd_sc_hd__dfrtp_1 _649_ (.CLK(clknet_2_0__leaf_clk),
    .D(\Adder.cla_16_bit.Sum[7] ),
    .RESET_B(_007_),
    .Q(net31));
 sky130_fd_sc_hd__dfrtp_1 _650_ (.CLK(clknet_2_0__leaf_clk),
    .D(\Adder.cla_16_bit.Sum[8] ),
    .RESET_B(_008_),
    .Q(net32));
 sky130_fd_sc_hd__dfrtp_1 _651_ (.CLK(clknet_2_1__leaf_clk),
    .D(\Adder.cla_16_bit.Sum[9] ),
    .RESET_B(_009_),
    .Q(net33));
 sky130_fd_sc_hd__dfrtp_1 _652_ (.CLK(clknet_2_2__leaf_clk),
    .D(\Adder.cla_16_bit.Sum[10] ),
    .RESET_B(_010_),
    .Q(net19));
 sky130_fd_sc_hd__dfrtp_1 _653_ (.CLK(clknet_2_1__leaf_clk),
    .D(\Adder.cla_16_bit.Sum[11] ),
    .RESET_B(_011_),
    .Q(net20));
 sky130_fd_sc_hd__dfrtp_1 _654_ (.CLK(clknet_2_1__leaf_clk),
    .D(\Adder.cla_16_bit.Sum[12] ),
    .RESET_B(_012_),
    .Q(net21));
 sky130_fd_sc_hd__dfrtp_1 _655_ (.CLK(clknet_2_1__leaf_clk),
    .D(\Adder.cla_16_bit.Sum[13] ),
    .RESET_B(_013_),
    .Q(net22));
 sky130_fd_sc_hd__dfrtp_1 _656_ (.CLK(clknet_2_1__leaf_clk),
    .D(\Adder.cla_16_bit.Sum[14] ),
    .RESET_B(_014_),
    .Q(net23));
 sky130_fd_sc_hd__dfrtp_1 _657_ (.CLK(clknet_2_1__leaf_clk),
    .D(\Adder.cla_16_bit.Sum[15] ),
    .RESET_B(_015_),
    .Q(net24));
 sky130_fd_sc_hd__dfrtp_4 _658_ (.CLK(clknet_2_1__leaf_clk),
    .D(net1),
    .RESET_B(_016_),
    .Q(\A_ff[0] ));
 sky130_fd_sc_hd__dfrtp_4 _659_ (.CLK(clknet_2_2__leaf_clk),
    .D(net2),
    .RESET_B(_017_),
    .Q(\A_ff[1] ));
 sky130_fd_sc_hd__dfrtp_4 _660_ (.CLK(clknet_2_1__leaf_clk),
    .D(net3),
    .RESET_B(_018_),
    .Q(\A_ff[2] ));
 sky130_fd_sc_hd__dfrtp_4 _661_ (.CLK(clknet_2_1__leaf_clk),
    .D(net4),
    .RESET_B(_019_),
    .Q(\A_ff[3] ));
 sky130_fd_sc_hd__dfrtp_4 _662_ (.CLK(clknet_2_1__leaf_clk),
    .D(net5),
    .RESET_B(_020_),
    .Q(\A_ff[4] ));
 sky130_fd_sc_hd__dfrtp_4 _663_ (.CLK(clknet_2_3__leaf_clk),
    .D(net6),
    .RESET_B(_021_),
    .Q(\A_ff[5] ));
 sky130_fd_sc_hd__dfrtp_4 _664_ (.CLK(clknet_2_2__leaf_clk),
    .D(net7),
    .RESET_B(_022_),
    .Q(\A_ff[6] ));
 sky130_fd_sc_hd__dfrtp_4 _665_ (.CLK(clknet_2_2__leaf_clk),
    .D(net8),
    .RESET_B(_023_),
    .Q(\A_ff[7] ));
 sky130_fd_sc_hd__dfrtp_4 _666_ (.CLK(clknet_2_2__leaf_clk),
    .D(net9),
    .RESET_B(_024_),
    .Q(\B_ff[0] ));
 sky130_fd_sc_hd__dfrtp_4 _667_ (.CLK(clknet_2_2__leaf_clk),
    .D(net10),
    .RESET_B(_025_),
    .Q(\B_ff[1] ));
 sky130_fd_sc_hd__dfrtp_4 _668_ (.CLK(clknet_2_3__leaf_clk),
    .D(net11),
    .RESET_B(_026_),
    .Q(\B_ff[2] ));
 sky130_fd_sc_hd__dfrtp_4 _669_ (.CLK(clknet_2_3__leaf_clk),
    .D(net12),
    .RESET_B(_027_),
    .Q(\B_ff[3] ));
 sky130_fd_sc_hd__dfrtp_2 _670_ (.CLK(clknet_2_3__leaf_clk),
    .D(net13),
    .RESET_B(_028_),
    .Q(\B_ff[4] ));
 sky130_fd_sc_hd__dfrtp_4 _671_ (.CLK(clknet_2_3__leaf_clk),
    .D(net14),
    .RESET_B(_029_),
    .Q(\B_ff[5] ));
 sky130_fd_sc_hd__dfrtp_1 _672_ (.CLK(clknet_2_3__leaf_clk),
    .D(net15),
    .RESET_B(_030_),
    .Q(\B_ff[6] ));
 sky130_fd_sc_hd__dfrtp_1 _673_ (.CLK(clknet_2_3__leaf_clk),
    .D(net16),
    .RESET_B(_031_),
    .Q(\B_ff[7] ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_155 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(A[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(A[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(A[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(A[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(A[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(A[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(A[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(A[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(B[0]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(B[1]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(B[2]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(B[3]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(B[4]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(B[5]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(B[6]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(B[7]),
    .X(net16));
 sky130_fd_sc_hd__buf_12 input17 (.A(reset),
    .X(net17));
 sky130_fd_sc_hd__buf_1 output18 (.A(net18),
    .X(Output[0]));
 sky130_fd_sc_hd__buf_1 output19 (.A(net19),
    .X(Output[10]));
 sky130_fd_sc_hd__buf_1 output20 (.A(net20),
    .X(Output[11]));
 sky130_fd_sc_hd__buf_1 output21 (.A(net21),
    .X(Output[12]));
 sky130_fd_sc_hd__buf_1 output22 (.A(net22),
    .X(Output[13]));
 sky130_fd_sc_hd__buf_1 output23 (.A(net23),
    .X(Output[14]));
 sky130_fd_sc_hd__buf_1 output24 (.A(net24),
    .X(Output[15]));
 sky130_fd_sc_hd__buf_1 output25 (.A(net25),
    .X(Output[1]));
 sky130_fd_sc_hd__buf_1 output26 (.A(net26),
    .X(Output[2]));
 sky130_fd_sc_hd__buf_1 output27 (.A(net27),
    .X(Output[3]));
 sky130_fd_sc_hd__buf_1 output28 (.A(net28),
    .X(Output[4]));
 sky130_fd_sc_hd__buf_1 output29 (.A(net29),
    .X(Output[5]));
 sky130_fd_sc_hd__buf_1 output30 (.A(net30),
    .X(Output[6]));
 sky130_fd_sc_hd__buf_1 output31 (.A(net31),
    .X(Output[7]));
 sky130_fd_sc_hd__buf_1 output32 (.A(net32),
    .X(Output[8]));
 sky130_fd_sc_hd__buf_1 output33 (.A(net33),
    .X(Output[9]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload0 (.A(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__bufinv_16 clkload1 (.A(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkinv_2 clkload2 (.A(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__decap_4 FILLER_0_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_172 ();
endmodule
