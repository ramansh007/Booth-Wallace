magic
tech sky130A
magscale 1 2
timestamp 1769689532
<< viali >>
rect 1685 18377 1719 18411
rect 2513 18377 2547 18411
rect 5825 18377 5859 18411
rect 1409 18241 1443 18275
rect 1869 18241 1903 18275
rect 2329 18241 2363 18275
rect 3433 18241 3467 18275
rect 4537 18241 4571 18275
rect 5641 18241 5675 18275
rect 6009 18241 6043 18275
rect 8677 18241 8711 18275
rect 8953 18241 8987 18275
rect 10241 18241 10275 18275
rect 11069 18241 11103 18275
rect 11161 18241 11195 18275
rect 12265 18241 12299 18275
rect 13553 18241 13587 18275
rect 14473 18241 14507 18275
rect 15761 18241 15795 18275
rect 16865 18241 16899 18275
rect 17509 18241 17543 18275
rect 6377 18173 6411 18207
rect 6653 18173 6687 18207
rect 8401 18173 8435 18207
rect 4721 18105 4755 18139
rect 1593 18037 1627 18071
rect 3617 18037 3651 18071
rect 6193 18037 6227 18071
rect 8493 18037 8527 18071
rect 9137 18037 9171 18071
rect 10057 18037 10091 18071
rect 10977 18037 11011 18071
rect 11345 18037 11379 18071
rect 12449 18037 12483 18071
rect 13369 18037 13403 18071
rect 14657 18037 14691 18071
rect 15577 18037 15611 18071
rect 16681 18037 16715 18071
rect 17325 18037 17359 18071
rect 9045 17765 9079 17799
rect 1409 17697 1443 17731
rect 4629 17697 4663 17731
rect 6745 17697 6779 17731
rect 7021 17697 7055 17731
rect 9781 17697 9815 17731
rect 10057 17697 10091 17731
rect 11897 17697 11931 17731
rect 14657 17697 14691 17731
rect 14933 17697 14967 17731
rect 3985 17629 4019 17663
rect 4537 17629 4571 17663
rect 9137 17629 9171 17663
rect 14289 17629 14323 17663
rect 16865 17629 16899 17663
rect 1685 17561 1719 17595
rect 3433 17561 3467 17595
rect 4905 17561 4939 17595
rect 6653 17561 6687 17595
rect 8769 17561 8803 17595
rect 11805 17561 11839 17595
rect 12173 17561 12207 17595
rect 13921 17561 13955 17595
rect 16681 17561 16715 17595
rect 3893 17493 3927 17527
rect 4445 17493 4479 17527
rect 14197 17493 14231 17527
rect 16957 17493 16991 17527
rect 1409 17289 1443 17323
rect 2237 17289 2271 17323
rect 3525 17289 3559 17323
rect 6469 17289 6503 17323
rect 7113 17289 7147 17323
rect 12541 17289 12575 17323
rect 15669 17289 15703 17323
rect 8217 17221 8251 17255
rect 1593 17153 1627 17187
rect 2145 17153 2179 17187
rect 6561 17153 6595 17187
rect 7021 17153 7055 17187
rect 10885 17153 10919 17187
rect 12449 17153 12483 17187
rect 13001 17153 13035 17187
rect 15577 17153 15611 17187
rect 4997 17085 5031 17119
rect 5273 17085 5307 17119
rect 7941 17085 7975 17119
rect 9965 17085 9999 17119
rect 13277 17085 13311 17119
rect 15025 17085 15059 17119
rect 10977 16949 11011 16983
rect 3433 16745 3467 16779
rect 9137 16745 9171 16779
rect 10130 16745 10164 16779
rect 15209 16677 15243 16711
rect 3157 16609 3191 16643
rect 9873 16609 9907 16643
rect 15761 16609 15795 16643
rect 16037 16609 16071 16643
rect 1593 16541 1627 16575
rect 3065 16541 3099 16575
rect 4077 16541 4111 16575
rect 4169 16541 4203 16575
rect 4261 16541 4295 16575
rect 4445 16541 4479 16575
rect 9229 16541 9263 16575
rect 13001 16541 13035 16575
rect 13277 16541 13311 16575
rect 14933 16541 14967 16575
rect 15117 16541 15151 16575
rect 15393 16541 15427 16575
rect 15577 16541 15611 16575
rect 11897 16473 11931 16507
rect 1409 16405 1443 16439
rect 3801 16405 3835 16439
rect 12817 16405 12851 16439
rect 13185 16405 13219 16439
rect 15025 16405 15059 16439
rect 17509 16405 17543 16439
rect 2881 16201 2915 16235
rect 5181 16201 5215 16235
rect 5825 16201 5859 16235
rect 8769 16201 8803 16235
rect 4353 16133 4387 16167
rect 7389 16133 7423 16167
rect 13369 16133 13403 16167
rect 14381 16133 14415 16167
rect 15025 16133 15059 16167
rect 1593 16065 1627 16099
rect 2145 16065 2179 16099
rect 5549 16065 5583 16099
rect 5825 16065 5859 16099
rect 6009 16065 6043 16099
rect 6377 16065 6411 16099
rect 6561 16065 6595 16099
rect 7021 16065 7055 16099
rect 7205 16065 7239 16099
rect 7297 16065 7331 16099
rect 7481 16065 7515 16099
rect 8677 16065 8711 16099
rect 8861 16065 8895 16099
rect 12265 16065 12299 16099
rect 12449 16065 12483 16099
rect 12633 16065 12667 16099
rect 12817 16065 12851 16099
rect 13277 16065 13311 16099
rect 13737 16065 13771 16099
rect 13921 16065 13955 16099
rect 14013 16065 14047 16099
rect 14197 16065 14231 16099
rect 14657 16065 14691 16099
rect 14841 16065 14875 16099
rect 14933 16065 14967 16099
rect 15117 16065 15151 16099
rect 15669 16065 15703 16099
rect 15853 16065 15887 16099
rect 16865 16065 16899 16099
rect 4629 15997 4663 16031
rect 5641 15997 5675 16031
rect 6745 15997 6779 16031
rect 6837 15997 6871 16031
rect 12541 15997 12575 16031
rect 13553 15997 13587 16031
rect 14473 15997 14507 16031
rect 15761 15997 15795 16031
rect 12909 15929 12943 15963
rect 1409 15861 1443 15895
rect 2237 15861 2271 15895
rect 12081 15861 12115 15895
rect 13737 15861 13771 15895
rect 16957 15861 16991 15895
rect 1409 15657 1443 15691
rect 3341 15657 3375 15691
rect 6653 15657 6687 15691
rect 9505 15657 9539 15691
rect 11529 15657 11563 15691
rect 13553 15657 13587 15691
rect 15025 15657 15059 15691
rect 15209 15589 15243 15623
rect 4261 15521 4295 15555
rect 7849 15521 7883 15555
rect 8033 15521 8067 15555
rect 8493 15521 8527 15555
rect 10793 15521 10827 15555
rect 11253 15521 11287 15555
rect 14473 15521 14507 15555
rect 15761 15521 15795 15555
rect 17233 15521 17267 15555
rect 3157 15453 3191 15487
rect 3525 15453 3559 15487
rect 3617 15453 3651 15487
rect 4169 15453 4203 15487
rect 4445 15453 4479 15487
rect 4720 15453 4754 15487
rect 4813 15453 4847 15487
rect 6193 15453 6227 15487
rect 6377 15453 6411 15487
rect 6469 15453 6503 15487
rect 7679 15453 7713 15487
rect 8401 15453 8435 15487
rect 9134 15453 9168 15487
rect 9597 15453 9631 15487
rect 9965 15453 9999 15487
rect 10057 15453 10091 15487
rect 10517 15453 10551 15487
rect 10701 15453 10735 15487
rect 11161 15453 11195 15487
rect 11437 15453 11471 15487
rect 11621 15453 11655 15487
rect 12173 15453 12207 15487
rect 12357 15453 12391 15487
rect 12449 15453 12483 15487
rect 12541 15453 12575 15487
rect 12725 15453 12759 15487
rect 12909 15453 12943 15487
rect 13001 15453 13035 15487
rect 13369 15453 13403 15487
rect 14197 15453 14231 15487
rect 14381 15453 14415 15487
rect 14657 15453 14691 15487
rect 14841 15453 14875 15487
rect 14933 15453 14967 15487
rect 15117 15453 15151 15487
rect 15209 15453 15243 15487
rect 15393 15453 15427 15487
rect 17509 15453 17543 15487
rect 2881 15385 2915 15419
rect 3341 15385 3375 15419
rect 6837 15385 6871 15419
rect 7021 15385 7055 15419
rect 9781 15385 9815 15419
rect 13185 15385 13219 15419
rect 13277 15385 13311 15419
rect 3801 15317 3835 15351
rect 7481 15317 7515 15351
rect 8953 15317 8987 15351
rect 9137 15317 9171 15351
rect 10425 15317 10459 15351
rect 10517 15317 10551 15351
rect 14289 15317 14323 15351
rect 1409 15113 1443 15147
rect 4261 15113 4295 15147
rect 8033 15113 8067 15147
rect 8493 15113 8527 15147
rect 8661 15113 8695 15147
rect 10701 15113 10735 15147
rect 12909 15113 12943 15147
rect 13921 15113 13955 15147
rect 16037 15113 16071 15147
rect 6929 15045 6963 15079
rect 7113 15045 7147 15079
rect 7573 15045 7607 15079
rect 8861 15045 8895 15079
rect 15025 15045 15059 15079
rect 4537 14977 4571 15011
rect 7481 14977 7515 15011
rect 7665 14977 7699 15011
rect 7849 14977 7883 15011
rect 8125 14977 8159 15011
rect 10149 14977 10183 15011
rect 10425 14977 10459 15011
rect 12173 14977 12207 15011
rect 12449 14977 12483 15011
rect 12633 14977 12667 15011
rect 12725 14977 12759 15011
rect 12909 14977 12943 15011
rect 13829 14977 13863 15011
rect 14105 14977 14139 15011
rect 14197 14977 14231 15011
rect 14381 14977 14415 15011
rect 14565 14977 14599 15011
rect 14749 14977 14783 15011
rect 14933 14977 14967 15011
rect 15301 14977 15335 15011
rect 15669 14977 15703 15011
rect 16681 14977 16715 15011
rect 2881 14909 2915 14943
rect 3157 14909 3191 14943
rect 4445 14909 4479 14943
rect 4629 14909 4663 14943
rect 4721 14909 4755 14943
rect 10241 14909 10275 14943
rect 10701 14909 10735 14943
rect 14657 14909 14691 14943
rect 15025 14909 15059 14943
rect 7849 14841 7883 14875
rect 11989 14841 12023 14875
rect 14105 14841 14139 14875
rect 16221 14841 16255 14875
rect 6745 14773 6779 14807
rect 8677 14773 8711 14807
rect 9781 14773 9815 14807
rect 10517 14773 10551 14807
rect 15209 14773 15243 14807
rect 16037 14773 16071 14807
rect 16773 14773 16807 14807
rect 2421 14569 2455 14603
rect 3985 14569 4019 14603
rect 4445 14569 4479 14603
rect 5641 14569 5675 14603
rect 9965 14569 9999 14603
rect 10885 14569 10919 14603
rect 11069 14569 11103 14603
rect 11437 14569 11471 14603
rect 4721 14501 4755 14535
rect 10517 14433 10551 14467
rect 1593 14365 1627 14399
rect 2513 14365 2547 14399
rect 3985 14365 4019 14399
rect 4169 14365 4203 14399
rect 4997 14365 5031 14399
rect 5365 14365 5399 14399
rect 5549 14365 5583 14399
rect 5641 14365 5675 14399
rect 5825 14365 5859 14399
rect 6101 14365 6135 14399
rect 6285 14365 6319 14399
rect 6377 14365 6411 14399
rect 6652 14365 6686 14399
rect 6745 14365 6779 14399
rect 9965 14365 9999 14399
rect 10149 14365 10183 14399
rect 10609 14365 10643 14399
rect 11069 14365 11103 14399
rect 11161 14365 11195 14399
rect 15669 14365 15703 14399
rect 4429 14297 4463 14331
rect 4629 14297 4663 14331
rect 4721 14297 4755 14331
rect 5457 14297 5491 14331
rect 5917 14297 5951 14331
rect 15945 14297 15979 14331
rect 1409 14229 1443 14263
rect 4261 14229 4295 14263
rect 4905 14229 4939 14263
rect 17417 14229 17451 14263
rect 1409 14025 1443 14059
rect 9781 14025 9815 14059
rect 11161 14025 11195 14059
rect 12265 14025 12299 14059
rect 12633 14025 12667 14059
rect 13461 14025 13495 14059
rect 14289 14025 14323 14059
rect 14565 14025 14599 14059
rect 16865 14025 16899 14059
rect 10057 13957 10091 13991
rect 12725 13957 12759 13991
rect 15025 13957 15059 13991
rect 15853 13957 15887 13991
rect 6745 13889 6779 13923
rect 9137 13889 9171 13923
rect 9689 13889 9723 13923
rect 9873 13889 9907 13923
rect 9965 13889 9999 13923
rect 10149 13889 10183 13923
rect 10609 13889 10643 13923
rect 11069 13889 11103 13923
rect 11253 13889 11287 13923
rect 13093 13889 13127 13923
rect 13369 13889 13403 13923
rect 14197 13889 14231 13923
rect 14473 13889 14507 13923
rect 14749 13889 14783 13923
rect 15209 13889 15243 13923
rect 15669 13889 15703 13923
rect 17049 13889 17083 13923
rect 2881 13821 2915 13855
rect 3157 13821 3191 13855
rect 6837 13821 6871 13855
rect 9321 13821 9355 13855
rect 9419 13821 9453 13855
rect 10701 13821 10735 13855
rect 12909 13821 12943 13855
rect 13185 13821 13219 13855
rect 16681 13821 16715 13855
rect 10241 13753 10275 13787
rect 6469 13685 6503 13719
rect 8953 13685 8987 13719
rect 14933 13685 14967 13719
rect 15393 13685 15427 13719
rect 15485 13685 15519 13719
rect 17233 13685 17267 13719
rect 2329 13481 2363 13515
rect 2973 13481 3007 13515
rect 5549 13481 5583 13515
rect 6377 13481 6411 13515
rect 8033 13481 8067 13515
rect 11161 13481 11195 13515
rect 6193 13413 6227 13447
rect 7941 13413 7975 13447
rect 14197 13413 14231 13447
rect 3341 13345 3375 13379
rect 4905 13345 4939 13379
rect 5365 13345 5399 13379
rect 7665 13345 7699 13379
rect 8493 13345 8527 13379
rect 11529 13345 11563 13379
rect 16405 13345 16439 13379
rect 1593 13277 1627 13311
rect 2421 13277 2455 13311
rect 3249 13277 3283 13311
rect 5180 13277 5214 13311
rect 5266 13277 5300 13311
rect 5641 13277 5675 13311
rect 6101 13277 6135 13311
rect 6285 13277 6319 13311
rect 6377 13277 6411 13311
rect 6561 13277 6595 13311
rect 7573 13277 7607 13311
rect 8401 13277 8435 13311
rect 8953 13277 8987 13311
rect 11345 13277 11379 13311
rect 11897 13277 11931 13311
rect 13553 13277 13587 13311
rect 14381 13277 14415 13311
rect 14749 13277 14783 13311
rect 14841 13277 14875 13311
rect 15393 13277 15427 13311
rect 15761 13277 15795 13311
rect 16221 13277 16255 13311
rect 16773 13277 16807 13311
rect 16865 13277 16899 13311
rect 11989 13209 12023 13243
rect 1409 13141 1443 13175
rect 5365 13141 5399 13175
rect 1409 12937 1443 12971
rect 3525 12937 3559 12971
rect 8309 12937 8343 12971
rect 10149 12937 10183 12971
rect 13461 12937 13495 12971
rect 14289 12937 14323 12971
rect 15209 12937 15243 12971
rect 16221 12937 16255 12971
rect 8125 12869 8159 12903
rect 8861 12869 8895 12903
rect 12081 12869 12115 12903
rect 14611 12869 14645 12903
rect 14749 12869 14783 12903
rect 14841 12869 14875 12903
rect 3157 12801 3191 12835
rect 3433 12801 3467 12835
rect 3617 12801 3651 12835
rect 4751 12801 4785 12835
rect 4905 12801 4939 12835
rect 5273 12801 5307 12835
rect 5365 12801 5399 12835
rect 5457 12801 5491 12835
rect 5641 12801 5675 12835
rect 8217 12801 8251 12835
rect 8493 12801 8527 12835
rect 11069 12801 11103 12835
rect 11989 12801 12023 12835
rect 12173 12801 12207 12835
rect 12265 12801 12299 12835
rect 12449 12801 12483 12835
rect 12541 12801 12575 12835
rect 12633 12801 12667 12835
rect 12817 12801 12851 12835
rect 13921 12801 13955 12835
rect 14473 12801 14507 12835
rect 14933 12801 14967 12835
rect 15577 12801 15611 12835
rect 16129 12801 16163 12835
rect 16405 12801 16439 12835
rect 16865 12801 16899 12835
rect 16957 12801 16991 12835
rect 2881 12733 2915 12767
rect 4997 12733 5031 12767
rect 11161 12733 11195 12767
rect 13001 12733 13035 12767
rect 13553 12733 13587 12767
rect 13645 12733 13679 12767
rect 14013 12733 14047 12767
rect 15485 12733 15519 12767
rect 17325 12733 17359 12767
rect 4537 12665 4571 12699
rect 8493 12665 8527 12699
rect 10701 12665 10735 12699
rect 13093 12665 13127 12699
rect 15117 12665 15151 12699
rect 6653 12597 6687 12631
rect 13921 12597 13955 12631
rect 15393 12597 15427 12631
rect 16681 12597 16715 12631
rect 2237 12393 2271 12427
rect 3157 12393 3191 12427
rect 4077 12393 4111 12427
rect 5917 12393 5951 12427
rect 7113 12393 7147 12427
rect 16405 12393 16439 12427
rect 6285 12325 6319 12359
rect 7297 12325 7331 12359
rect 4721 12257 4755 12291
rect 6929 12257 6963 12291
rect 17049 12257 17083 12291
rect 1593 12189 1627 12223
rect 2145 12189 2179 12223
rect 3341 12189 3375 12223
rect 3617 12189 3651 12223
rect 4261 12189 4295 12223
rect 4353 12189 4387 12223
rect 5917 12189 5951 12223
rect 6101 12189 6135 12223
rect 6193 12189 6227 12223
rect 6377 12189 6411 12223
rect 6837 12189 6871 12223
rect 16405 12189 16439 12223
rect 16589 12189 16623 12223
rect 16865 12189 16899 12223
rect 7573 12121 7607 12155
rect 1409 12053 1443 12087
rect 3525 12053 3559 12087
rect 6469 12053 6503 12087
rect 16681 12053 16715 12087
rect 3617 11849 3651 11883
rect 3709 11849 3743 11883
rect 7021 11849 7055 11883
rect 8033 11849 8067 11883
rect 10793 11849 10827 11883
rect 14381 11849 14415 11883
rect 14657 11849 14691 11883
rect 16129 11849 16163 11883
rect 4445 11781 4479 11815
rect 4721 11781 4755 11815
rect 8585 11781 8619 11815
rect 10149 11781 10183 11815
rect 11529 11781 11563 11815
rect 13185 11781 13219 11815
rect 13921 11781 13955 11815
rect 3341 11713 3375 11747
rect 3801 11713 3835 11747
rect 3893 11713 3927 11747
rect 4077 11713 4111 11747
rect 4169 11713 4203 11747
rect 4353 11713 4387 11747
rect 4537 11713 4571 11747
rect 4629 11713 4663 11747
rect 6929 11713 6963 11747
rect 7113 11713 7147 11747
rect 8217 11713 8251 11747
rect 8401 11713 8435 11747
rect 8493 11713 8527 11747
rect 8769 11713 8803 11747
rect 9045 11713 9079 11747
rect 9229 11713 9263 11747
rect 10333 11713 10367 11747
rect 10425 11713 10459 11747
rect 11161 11713 11195 11747
rect 11713 11713 11747 11747
rect 11989 11713 12023 11747
rect 12449 11713 12483 11747
rect 12725 11713 12759 11747
rect 12817 11713 12851 11747
rect 13001 11713 13035 11747
rect 13093 11713 13127 11747
rect 13277 11713 13311 11747
rect 14013 11713 14047 11747
rect 14654 11713 14688 11747
rect 15209 11713 15243 11747
rect 15393 11713 15427 11747
rect 15485 11713 15519 11747
rect 15669 11713 15703 11747
rect 15761 11713 15795 11747
rect 15853 11713 15887 11747
rect 16313 11713 16347 11747
rect 16497 11713 16531 11747
rect 16865 11713 16899 11747
rect 17141 11713 17175 11747
rect 17325 11713 17359 11747
rect 11253 11645 11287 11679
rect 12633 11645 12667 11679
rect 13737 11645 13771 11679
rect 15117 11645 15151 11679
rect 16129 11645 16163 11679
rect 10149 11577 10183 11611
rect 14473 11577 14507 11611
rect 11897 11509 11931 11543
rect 12265 11509 12299 11543
rect 15025 11509 15059 11543
rect 15945 11509 15979 11543
rect 16405 11509 16439 11543
rect 16681 11509 16715 11543
rect 1409 11305 1443 11339
rect 4813 11305 4847 11339
rect 5457 11305 5491 11339
rect 10793 11305 10827 11339
rect 15669 11305 15703 11339
rect 3801 11237 3835 11271
rect 8953 11237 8987 11271
rect 2881 11169 2915 11203
rect 3157 11169 3191 11203
rect 4261 11169 4295 11203
rect 5181 11169 5215 11203
rect 6653 11169 6687 11203
rect 7113 11169 7147 11203
rect 8493 11169 8527 11203
rect 8769 11169 8803 11203
rect 9229 11169 9263 11203
rect 10517 11169 10551 11203
rect 12633 11169 12667 11203
rect 13001 11169 13035 11203
rect 13369 11169 13403 11203
rect 15117 11169 15151 11203
rect 15853 11169 15887 11203
rect 3433 11101 3467 11135
rect 4169 11101 4203 11135
rect 5089 11101 5123 11135
rect 5365 11101 5399 11135
rect 5549 11101 5583 11135
rect 7021 11101 7055 11135
rect 8401 11101 8435 11135
rect 9321 11101 9355 11135
rect 10425 11101 10459 11135
rect 12541 11101 12575 11135
rect 13553 11101 13587 11135
rect 13921 11101 13955 11135
rect 14749 11101 14783 11135
rect 14933 11101 14967 11135
rect 15209 11101 15243 11135
rect 15301 11101 15335 11135
rect 15485 11101 15519 11135
rect 15577 11101 15611 11135
rect 16497 11101 16531 11135
rect 3341 11033 3375 11067
rect 12357 11033 12391 11067
rect 15853 11033 15887 11067
rect 16129 11033 16163 11067
rect 16313 11033 16347 11067
rect 13553 10965 13587 10999
rect 1409 10761 1443 10795
rect 15209 10761 15243 10795
rect 11253 10693 11287 10727
rect 1593 10625 1627 10659
rect 6377 10625 6411 10659
rect 11713 10625 11747 10659
rect 11897 10625 11931 10659
rect 15117 10625 15151 10659
rect 15301 10625 15335 10659
rect 16681 10625 16715 10659
rect 16773 10625 16807 10659
rect 6653 10557 6687 10591
rect 8401 10557 8435 10591
rect 16957 10557 16991 10591
rect 9781 10421 9815 10455
rect 11529 10421 11563 10455
rect 16865 10421 16899 10455
rect 1409 10217 1443 10251
rect 6653 10217 6687 10251
rect 15025 10217 15059 10251
rect 16405 10217 16439 10251
rect 3893 10149 3927 10183
rect 10517 10149 10551 10183
rect 14565 10149 14599 10183
rect 16681 10149 16715 10183
rect 2881 10081 2915 10115
rect 3801 10081 3835 10115
rect 10241 10081 10275 10115
rect 10701 10081 10735 10115
rect 15209 10081 15243 10115
rect 3157 10013 3191 10047
rect 6561 10013 6595 10047
rect 9965 10013 9999 10047
rect 10057 10013 10091 10047
rect 10517 10013 10551 10047
rect 10885 10013 10919 10047
rect 12357 10013 12391 10047
rect 12541 10013 12575 10047
rect 12633 10013 12667 10047
rect 12817 10013 12851 10047
rect 12909 10013 12943 10047
rect 13093 10013 13127 10047
rect 14565 10013 14599 10047
rect 14841 10013 14875 10047
rect 14933 10013 14967 10047
rect 16221 10013 16255 10047
rect 16313 10013 16347 10047
rect 16957 10013 16991 10047
rect 17049 10013 17083 10047
rect 17233 10013 17267 10047
rect 4261 9945 4295 9979
rect 16681 9945 16715 9979
rect 12449 9877 12483 9911
rect 12725 9877 12759 9911
rect 12909 9877 12943 9911
rect 14749 9877 14783 9911
rect 15209 9877 15243 9911
rect 16589 9877 16623 9911
rect 16865 9877 16899 9911
rect 17141 9877 17175 9911
rect 3249 9673 3283 9707
rect 4537 9673 4571 9707
rect 5089 9673 5123 9707
rect 10149 9673 10183 9707
rect 2421 9605 2455 9639
rect 3617 9605 3651 9639
rect 5257 9605 5291 9639
rect 5457 9605 5491 9639
rect 8125 9605 8159 9639
rect 13737 9605 13771 9639
rect 1593 9537 1627 9571
rect 2513 9537 2547 9571
rect 3433 9537 3467 9571
rect 3525 9537 3559 9571
rect 3801 9537 3835 9571
rect 4077 9537 4111 9571
rect 4353 9537 4387 9571
rect 4721 9537 4755 9571
rect 4905 9537 4939 9571
rect 4997 9537 5031 9571
rect 5825 9537 5859 9571
rect 6377 9537 6411 9571
rect 8769 9537 8803 9571
rect 9229 9537 9263 9571
rect 9781 9537 9815 9571
rect 10609 9537 10643 9571
rect 11713 9537 11747 9571
rect 11805 9537 11839 9571
rect 12265 9537 12299 9571
rect 12357 9537 12391 9571
rect 12541 9537 12575 9571
rect 12633 9537 12667 9571
rect 12909 9537 12943 9571
rect 13093 9537 13127 9571
rect 13461 9537 13495 9571
rect 13921 9537 13955 9571
rect 14013 9537 14047 9571
rect 14289 9537 14323 9571
rect 14565 9537 14599 9571
rect 14749 9537 14783 9571
rect 15025 9537 15059 9571
rect 15389 9543 15423 9577
rect 15577 9537 15611 9571
rect 15669 9537 15703 9571
rect 15761 9537 15795 9571
rect 15853 9537 15887 9571
rect 16681 9537 16715 9571
rect 16865 9537 16899 9571
rect 17049 9537 17083 9571
rect 17233 9537 17267 9571
rect 3893 9469 3927 9503
rect 4169 9469 4203 9503
rect 4261 9469 4295 9503
rect 8677 9469 8711 9503
rect 9505 9469 9539 9503
rect 9873 9469 9907 9503
rect 10517 9469 10551 9503
rect 11989 9469 12023 9503
rect 13185 9469 13219 9503
rect 13277 9469 13311 9503
rect 13645 9469 13679 9503
rect 13737 9469 13771 9503
rect 14473 9469 14507 9503
rect 15209 9469 15243 9503
rect 15301 9469 15335 9503
rect 16957 9469 16991 9503
rect 1409 9401 1443 9435
rect 14105 9401 14139 9435
rect 14381 9401 14415 9435
rect 5273 9333 5307 9367
rect 8493 9333 8527 9367
rect 9045 9333 9079 9367
rect 9413 9333 9447 9367
rect 10333 9333 10367 9367
rect 11897 9333 11931 9367
rect 12081 9333 12115 9367
rect 14841 9333 14875 9367
rect 17417 9333 17451 9367
rect 1409 9129 1443 9163
rect 4353 9129 4387 9163
rect 7113 9129 7147 9163
rect 8309 9129 8343 9163
rect 8677 9129 8711 9163
rect 12633 9129 12667 9163
rect 14381 9129 14415 9163
rect 15117 9129 15151 9163
rect 3801 9061 3835 9095
rect 4629 9061 4663 9095
rect 3157 8993 3191 9027
rect 6469 8993 6503 9027
rect 6745 8993 6779 9027
rect 8033 8993 8067 9027
rect 16589 8993 16623 9027
rect 16681 8993 16715 9027
rect 17049 8993 17083 9027
rect 4169 8925 4203 8959
rect 4537 8925 4571 8959
rect 4813 8925 4847 8959
rect 5549 8925 5583 8959
rect 6009 8925 6043 8959
rect 6837 8925 6871 8959
rect 7113 8925 7147 8959
rect 7297 8925 7331 8959
rect 7941 8925 7975 8959
rect 8401 8925 8435 8959
rect 8677 8925 8711 8959
rect 12357 8925 12391 8959
rect 12633 8925 12667 8959
rect 14289 8925 14323 8959
rect 14749 8925 14783 8959
rect 15025 8925 15059 8959
rect 15117 8925 15151 8959
rect 15301 8925 15335 8959
rect 17141 8925 17175 8959
rect 2881 8857 2915 8891
rect 4077 8857 4111 8891
rect 4721 8857 4755 8891
rect 8493 8857 8527 8891
rect 14841 8857 14875 8891
rect 17233 8857 17267 8891
rect 3985 8789 4019 8823
rect 5181 8789 5215 8823
rect 12449 8789 12483 8823
rect 14926 8789 14960 8823
rect 16405 8789 16439 8823
rect 1409 8585 1443 8619
rect 2237 8585 2271 8619
rect 5457 8585 5491 8619
rect 5733 8585 5767 8619
rect 9229 8585 9263 8619
rect 12081 8585 12115 8619
rect 12173 8517 12207 8551
rect 1593 8449 1627 8483
rect 2145 8449 2179 8483
rect 3249 8449 3283 8483
rect 5200 8449 5234 8483
rect 5365 8449 5399 8483
rect 5641 8449 5675 8483
rect 5733 8449 5767 8483
rect 5917 8449 5951 8483
rect 7205 8449 7239 8483
rect 7481 8449 7515 8483
rect 7665 8449 7699 8483
rect 7757 8449 7791 8483
rect 9413 8449 9447 8483
rect 9597 8449 9631 8483
rect 9689 8449 9723 8483
rect 12541 8449 12575 8483
rect 2881 8381 2915 8415
rect 3341 8381 3375 8415
rect 7297 8381 7331 8415
rect 12081 8381 12115 8415
rect 6837 8313 6871 8347
rect 7481 8313 7515 8347
rect 11621 8313 11655 8347
rect 12449 8245 12483 8279
rect 1409 8041 1443 8075
rect 7297 8041 7331 8075
rect 9965 8041 9999 8075
rect 16681 8041 16715 8075
rect 5549 7973 5583 8007
rect 7205 7973 7239 8007
rect 7389 7973 7423 8007
rect 7849 7973 7883 8007
rect 10057 7973 10091 8007
rect 16865 7973 16899 8007
rect 3157 7905 3191 7939
rect 5273 7905 5307 7939
rect 6929 7905 6963 7939
rect 9781 7905 9815 7939
rect 11069 7905 11103 7939
rect 11345 7905 11379 7939
rect 13093 7905 13127 7939
rect 16773 7905 16807 7939
rect 5181 7837 5215 7871
rect 6837 7837 6871 7871
rect 8124 7837 8158 7871
rect 8217 7837 8251 7871
rect 9689 7837 9723 7871
rect 14841 7837 14875 7871
rect 15761 7837 15795 7871
rect 15915 7837 15949 7871
rect 16129 7837 16163 7871
rect 16221 7837 16255 7871
rect 16497 7837 16531 7871
rect 2881 7769 2915 7803
rect 7757 7769 7791 7803
rect 10425 7769 10459 7803
rect 14657 7769 14691 7803
rect 17233 7769 17267 7803
rect 9321 7701 9355 7735
rect 14473 7701 14507 7735
rect 16313 7701 16347 7735
rect 1409 7497 1443 7531
rect 2329 7497 2363 7531
rect 9505 7497 9539 7531
rect 9597 7497 9631 7531
rect 10149 7497 10183 7531
rect 15577 7497 15611 7531
rect 12449 7429 12483 7463
rect 1593 7361 1627 7395
rect 2421 7361 2455 7395
rect 3801 7361 3835 7395
rect 4445 7361 4479 7395
rect 4721 7361 4755 7395
rect 4905 7361 4939 7395
rect 9137 7361 9171 7395
rect 9781 7361 9815 7395
rect 9965 7361 9999 7395
rect 10057 7361 10091 7395
rect 10241 7361 10275 7395
rect 12173 7361 12207 7395
rect 14565 7361 14599 7395
rect 15209 7361 15243 7395
rect 16865 7361 16899 7395
rect 3433 7293 3467 7327
rect 3709 7293 3743 7327
rect 4077 7293 4111 7327
rect 4537 7293 4571 7327
rect 9229 7293 9263 7327
rect 10885 7293 10919 7327
rect 14197 7293 14231 7327
rect 14657 7293 14691 7327
rect 14933 7293 14967 7327
rect 15117 7293 15151 7327
rect 16773 7293 16807 7327
rect 11161 7225 11195 7259
rect 4721 7157 4755 7191
rect 9965 7157 9999 7191
rect 11345 7157 11379 7191
rect 17233 7157 17267 7191
rect 1409 6953 1443 6987
rect 11069 6953 11103 6987
rect 13737 6953 13771 6987
rect 3157 6817 3191 6851
rect 4261 6817 4295 6851
rect 9321 6817 9355 6851
rect 11713 6817 11747 6851
rect 13369 6817 13403 6851
rect 13645 6817 13679 6851
rect 14381 6817 14415 6851
rect 16405 6817 16439 6851
rect 17233 6817 17267 6851
rect 3801 6749 3835 6783
rect 3893 6749 3927 6783
rect 4077 6749 4111 6783
rect 7389 6749 7423 6783
rect 7665 6749 7699 6783
rect 9229 6749 9263 6783
rect 9413 6749 9447 6783
rect 11529 6749 11563 6783
rect 11897 6749 11931 6783
rect 12081 6749 12115 6783
rect 13461 6749 13495 6783
rect 13829 6749 13863 6783
rect 13921 6749 13955 6783
rect 14565 6749 14599 6783
rect 14749 6749 14783 6783
rect 14841 6749 14875 6783
rect 15117 6749 15151 6783
rect 15209 6749 15243 6783
rect 17049 6749 17083 6783
rect 2881 6681 2915 6715
rect 7573 6681 7607 6715
rect 11437 6681 11471 6715
rect 12265 6681 12299 6715
rect 14933 6613 14967 6647
rect 1409 6409 1443 6443
rect 2329 6409 2363 6443
rect 4721 6409 4755 6443
rect 5825 6409 5859 6443
rect 9137 6409 9171 6443
rect 8677 6341 8711 6375
rect 12725 6341 12759 6375
rect 1593 6273 1627 6307
rect 2421 6273 2455 6307
rect 3985 6273 4019 6307
rect 4261 6273 4295 6307
rect 4353 6273 4387 6307
rect 4537 6273 4571 6307
rect 6100 6273 6134 6307
rect 6193 6273 6227 6307
rect 6745 6273 6779 6307
rect 7941 6273 7975 6307
rect 8125 6273 8159 6307
rect 8769 6273 8803 6307
rect 9873 6273 9907 6307
rect 11989 6273 12023 6307
rect 12636 6273 12670 6307
rect 12909 6273 12943 6307
rect 14473 6273 14507 6307
rect 14657 6273 14691 6307
rect 14749 6273 14783 6307
rect 3617 6205 3651 6239
rect 4077 6205 4111 6239
rect 6837 6205 6871 6239
rect 8585 6205 8619 6239
rect 10149 6205 10183 6239
rect 11805 6205 11839 6239
rect 11897 6205 11931 6239
rect 12357 6137 12391 6171
rect 6469 6069 6503 6103
rect 8033 6069 8067 6103
rect 9965 6069 9999 6103
rect 10057 6069 10091 6103
rect 12909 6069 12943 6103
rect 14473 6069 14507 6103
rect 4261 5865 4295 5899
rect 5641 5865 5675 5899
rect 6193 5865 6227 5899
rect 7665 5865 7699 5899
rect 9597 5865 9631 5899
rect 10333 5865 10367 5899
rect 10517 5865 10551 5899
rect 11161 5865 11195 5899
rect 12449 5865 12483 5899
rect 13093 5865 13127 5899
rect 16221 5865 16255 5899
rect 16497 5865 16531 5899
rect 6377 5797 6411 5831
rect 9505 5797 9539 5831
rect 14933 5797 14967 5831
rect 6009 5729 6043 5763
rect 11621 5729 11655 5763
rect 11713 5729 11747 5763
rect 12284 5729 12318 5763
rect 12909 5729 12943 5763
rect 13553 5729 13587 5763
rect 13737 5729 13771 5763
rect 14749 5729 14783 5763
rect 15577 5729 15611 5763
rect 16129 5729 16163 5763
rect 16681 5729 16715 5763
rect 1593 5661 1627 5695
rect 4445 5661 4479 5695
rect 4721 5661 4755 5695
rect 5917 5661 5951 5695
rect 7481 5661 7515 5695
rect 7635 5661 7669 5695
rect 7941 5661 7975 5695
rect 8125 5661 8159 5695
rect 8217 5661 8251 5695
rect 8309 5661 8343 5695
rect 8493 5661 8527 5695
rect 9229 5661 9263 5695
rect 9321 5661 9355 5695
rect 9781 5661 9815 5695
rect 9873 5661 9907 5695
rect 12081 5661 12115 5695
rect 12633 5661 12667 5695
rect 12725 5661 12759 5695
rect 13001 5661 13035 5695
rect 14565 5661 14599 5695
rect 15393 5661 15427 5695
rect 15945 5661 15979 5695
rect 16773 5661 16807 5695
rect 6653 5593 6687 5627
rect 9505 5593 9539 5627
rect 10701 5593 10735 5627
rect 12173 5593 12207 5627
rect 12357 5593 12391 5627
rect 13461 5593 13495 5627
rect 14473 5593 14507 5627
rect 15301 5593 15335 5627
rect 16313 5593 16347 5627
rect 1409 5525 1443 5559
rect 4629 5525 4663 5559
rect 8677 5525 8711 5559
rect 10241 5525 10275 5559
rect 10501 5525 10535 5559
rect 11529 5525 11563 5559
rect 14105 5525 14139 5559
rect 1409 5321 1443 5355
rect 5365 5321 5399 5355
rect 7757 5321 7791 5355
rect 8125 5321 8159 5355
rect 10977 5321 11011 5355
rect 12541 5321 12575 5355
rect 16405 5321 16439 5355
rect 5701 5253 5735 5287
rect 5917 5253 5951 5287
rect 7573 5253 7607 5287
rect 3157 5185 3191 5219
rect 3893 5185 3927 5219
rect 4628 5185 4662 5219
rect 4721 5185 4755 5219
rect 5181 5185 5215 5219
rect 5457 5185 5491 5219
rect 7205 5185 7239 5219
rect 8585 5185 8619 5219
rect 8769 5185 8803 5219
rect 10241 5185 10275 5219
rect 10425 5185 10459 5219
rect 10609 5185 10643 5219
rect 10701 5185 10735 5219
rect 10793 5185 10827 5219
rect 12725 5185 12759 5219
rect 12817 5185 12851 5219
rect 13093 5185 13127 5219
rect 14289 5185 14323 5219
rect 14381 5185 14415 5219
rect 14657 5185 14691 5219
rect 15289 5185 15323 5219
rect 15485 5185 15519 5219
rect 16037 5185 16071 5219
rect 16681 5185 16715 5219
rect 16865 5185 16899 5219
rect 2881 5117 2915 5151
rect 3985 5117 4019 5151
rect 4353 5117 4387 5151
rect 4997 5117 5031 5151
rect 7389 5117 7423 5151
rect 8217 5117 8251 5151
rect 8401 5117 8435 5151
rect 15393 5117 15427 5151
rect 16129 5117 16163 5151
rect 3525 5049 3559 5083
rect 5549 5049 5583 5083
rect 7205 5049 7239 5083
rect 10057 5049 10091 5083
rect 14105 5049 14139 5083
rect 5733 4981 5767 5015
rect 8677 4981 8711 5015
rect 10241 4981 10275 5015
rect 13001 4981 13035 5015
rect 14565 4981 14599 5015
rect 16037 4981 16071 5015
rect 16681 4981 16715 5015
rect 2329 4777 2363 4811
rect 10885 4777 10919 4811
rect 11253 4777 11287 4811
rect 16773 4777 16807 4811
rect 9689 4709 9723 4743
rect 16681 4709 16715 4743
rect 16865 4709 16899 4743
rect 9321 4641 9355 4675
rect 10149 4641 10183 4675
rect 10609 4641 10643 4675
rect 10793 4641 10827 4675
rect 11161 4641 11195 4675
rect 16221 4641 16255 4675
rect 1593 4573 1627 4607
rect 2421 4573 2455 4607
rect 6193 4573 6227 4607
rect 6377 4573 6411 4607
rect 8953 4573 8987 4607
rect 9137 4573 9171 4607
rect 9229 4573 9263 4607
rect 9505 4573 9539 4607
rect 10517 4573 10551 4607
rect 11253 4573 11287 4607
rect 16313 4573 16347 4607
rect 17233 4573 17267 4607
rect 1409 4437 1443 4471
rect 6193 4437 6227 4471
rect 4353 4233 4387 4267
rect 8677 4233 8711 4267
rect 11069 4233 11103 4267
rect 12725 4233 12759 4267
rect 13461 4233 13495 4267
rect 14841 4233 14875 4267
rect 3341 4165 3375 4199
rect 5917 4165 5951 4199
rect 7113 4165 7147 4199
rect 13369 4165 13403 4199
rect 3157 4097 3191 4131
rect 3433 4097 3467 4131
rect 4077 4097 4111 4131
rect 6101 4097 6135 4131
rect 6193 4097 6227 4131
rect 6745 4097 6779 4131
rect 7021 4097 7055 4131
rect 7205 4097 7239 4131
rect 8309 4097 8343 4131
rect 8401 4097 8435 4131
rect 8493 4097 8527 4131
rect 12265 4097 12299 4131
rect 12403 4097 12437 4131
rect 12633 4097 12667 4131
rect 13001 4097 13035 4131
rect 13277 4097 13311 4131
rect 13737 4097 13771 4131
rect 13829 4097 13863 4131
rect 14782 4097 14816 4131
rect 15577 4097 15611 4131
rect 15669 4097 15703 4131
rect 1409 4029 1443 4063
rect 2881 4029 2915 4063
rect 4169 4029 4203 4063
rect 4813 4029 4847 4063
rect 6837 4029 6871 4063
rect 12081 4029 12115 4063
rect 12909 4029 12943 4063
rect 13645 4029 13679 4063
rect 15301 4029 15335 4063
rect 15393 4029 15427 4063
rect 3709 3961 3743 3995
rect 4537 3961 4571 3995
rect 5917 3961 5951 3995
rect 10701 3961 10735 3995
rect 14657 3961 14691 3995
rect 6469 3893 6503 3927
rect 11069 3893 11103 3927
rect 11253 3893 11287 3927
rect 12541 3893 12575 3927
rect 15209 3893 15243 3927
rect 15485 3893 15519 3927
rect 5917 3689 5951 3723
rect 8309 3689 8343 3723
rect 8493 3689 8527 3723
rect 10701 3689 10735 3723
rect 13001 3689 13035 3723
rect 13369 3689 13403 3723
rect 13737 3689 13771 3723
rect 13829 3689 13863 3723
rect 14841 3689 14875 3723
rect 15577 3689 15611 3723
rect 7849 3621 7883 3655
rect 15025 3621 15059 3655
rect 16037 3621 16071 3655
rect 3433 3553 3467 3587
rect 6377 3553 6411 3587
rect 9229 3553 9263 3587
rect 9321 3553 9355 3587
rect 11161 3553 11195 3587
rect 12265 3553 12299 3587
rect 13921 3553 13955 3587
rect 14381 3553 14415 3587
rect 14933 3553 14967 3587
rect 1593 3485 1627 3519
rect 3249 3485 3283 3519
rect 6285 3485 6319 3519
rect 7481 3485 7515 3519
rect 7665 3485 7699 3519
rect 8124 3485 8158 3519
rect 8217 3485 8251 3519
rect 9137 3485 9171 3519
rect 9413 3485 9447 3519
rect 10609 3485 10643 3519
rect 11069 3485 11103 3519
rect 11437 3485 11471 3519
rect 11621 3485 11655 3519
rect 12449 3485 12483 3519
rect 12725 3485 12759 3519
rect 12909 3485 12943 3519
rect 13185 3485 13219 3519
rect 13461 3485 13495 3519
rect 13645 3485 13679 3519
rect 14289 3485 14323 3519
rect 14565 3485 14599 3519
rect 14657 3485 14691 3519
rect 15452 3485 15486 3519
rect 15853 3485 15887 3519
rect 7573 3417 7607 3451
rect 8461 3417 8495 3451
rect 8677 3417 8711 3451
rect 15669 3417 15703 3451
rect 1409 3349 1443 3383
rect 3065 3349 3099 3383
rect 8953 3349 8987 3383
rect 15393 3349 15427 3383
rect 9866 3145 9900 3179
rect 10609 3145 10643 3179
rect 11713 3145 11747 3179
rect 12449 3145 12483 3179
rect 15117 3145 15151 3179
rect 3893 3077 3927 3111
rect 9781 3077 9815 3111
rect 1593 3009 1627 3043
rect 2145 3009 2179 3043
rect 4169 3009 4203 3043
rect 6009 3009 6043 3043
rect 7113 3009 7147 3043
rect 7389 3009 7423 3043
rect 7573 3009 7607 3043
rect 8585 3009 8619 3043
rect 9045 3009 9079 3043
rect 9229 3009 9263 3043
rect 9321 3009 9355 3043
rect 9689 3009 9723 3043
rect 9965 3009 9999 3043
rect 10057 3009 10091 3043
rect 10149 3009 10183 3043
rect 10793 3009 10827 3043
rect 10977 3009 11011 3043
rect 11253 3009 11287 3043
rect 11805 3009 11839 3043
rect 11989 3009 12023 3043
rect 13001 3009 13035 3043
rect 13645 3009 13679 3043
rect 14197 3009 14231 3043
rect 15301 3009 15335 3043
rect 15393 3009 15427 3043
rect 15669 3009 15703 3043
rect 2421 2941 2455 2975
rect 4261 2941 4295 2975
rect 5733 2941 5767 2975
rect 6745 2941 6779 2975
rect 7205 2941 7239 2975
rect 7481 2941 7515 2975
rect 8677 2941 8711 2975
rect 8861 2941 8895 2975
rect 10517 2941 10551 2975
rect 11529 2941 11563 2975
rect 12725 2941 12759 2975
rect 8217 2873 8251 2907
rect 10333 2873 10367 2907
rect 14381 2873 14415 2907
rect 15577 2873 15611 2907
rect 1409 2805 1443 2839
rect 2237 2805 2271 2839
rect 10793 2805 10827 2839
rect 12817 2805 12851 2839
rect 1409 2601 1443 2635
rect 3893 2601 3927 2635
rect 5365 2601 5399 2635
rect 11069 2601 11103 2635
rect 13185 2601 13219 2635
rect 3157 2465 3191 2499
rect 9965 2465 9999 2499
rect 3985 2397 4019 2431
rect 5273 2397 5307 2431
rect 9505 2397 9539 2431
rect 11161 2397 11195 2431
rect 13093 2397 13127 2431
rect 13277 2397 13311 2431
rect 2881 2329 2915 2363
<< metal1 >>
rect 1104 18522 17848 18544
rect 1104 18470 2658 18522
rect 2710 18470 2722 18522
rect 2774 18470 2786 18522
rect 2838 18470 2850 18522
rect 2902 18470 2914 18522
rect 2966 18470 2978 18522
rect 3030 18470 8658 18522
rect 8710 18470 8722 18522
rect 8774 18470 8786 18522
rect 8838 18470 8850 18522
rect 8902 18470 8914 18522
rect 8966 18470 8978 18522
rect 9030 18470 14658 18522
rect 14710 18470 14722 18522
rect 14774 18470 14786 18522
rect 14838 18470 14850 18522
rect 14902 18470 14914 18522
rect 14966 18470 14978 18522
rect 15030 18470 17848 18522
rect 1104 18448 17848 18470
rect 1210 18368 1216 18420
rect 1268 18408 1274 18420
rect 1673 18411 1731 18417
rect 1673 18408 1685 18411
rect 1268 18380 1685 18408
rect 1268 18368 1274 18380
rect 1673 18377 1685 18380
rect 1719 18377 1731 18411
rect 1673 18371 1731 18377
rect 2501 18411 2559 18417
rect 2501 18377 2513 18411
rect 2547 18408 2559 18411
rect 5718 18408 5724 18420
rect 2547 18380 5724 18408
rect 2547 18377 2559 18380
rect 2501 18371 2559 18377
rect 5718 18368 5724 18380
rect 5776 18368 5782 18420
rect 5813 18411 5871 18417
rect 5813 18377 5825 18411
rect 5859 18408 5871 18411
rect 7006 18408 7012 18420
rect 5859 18380 7012 18408
rect 5859 18377 5871 18380
rect 5813 18371 5871 18377
rect 7006 18368 7012 18380
rect 7064 18368 7070 18420
rect 6638 18340 6644 18352
rect 6012 18312 6644 18340
rect 1118 18232 1124 18284
rect 1176 18272 1182 18284
rect 1397 18275 1455 18281
rect 1397 18272 1409 18275
rect 1176 18244 1409 18272
rect 1176 18232 1182 18244
rect 1397 18241 1409 18244
rect 1443 18241 1455 18275
rect 1397 18235 1455 18241
rect 1857 18275 1915 18281
rect 1857 18241 1869 18275
rect 1903 18241 1915 18275
rect 1857 18235 1915 18241
rect 1872 18204 1900 18235
rect 2222 18232 2228 18284
rect 2280 18272 2286 18284
rect 2317 18275 2375 18281
rect 2317 18272 2329 18275
rect 2280 18244 2329 18272
rect 2280 18232 2286 18244
rect 2317 18241 2329 18244
rect 2363 18241 2375 18275
rect 2317 18235 2375 18241
rect 3326 18232 3332 18284
rect 3384 18272 3390 18284
rect 3421 18275 3479 18281
rect 3421 18272 3433 18275
rect 3384 18244 3433 18272
rect 3384 18232 3390 18244
rect 3421 18241 3433 18244
rect 3467 18241 3479 18275
rect 3421 18235 3479 18241
rect 4430 18232 4436 18284
rect 4488 18272 4494 18284
rect 4525 18275 4583 18281
rect 4525 18272 4537 18275
rect 4488 18244 4537 18272
rect 4488 18232 4494 18244
rect 4525 18241 4537 18244
rect 4571 18241 4583 18275
rect 4525 18235 4583 18241
rect 5534 18232 5540 18284
rect 5592 18272 5598 18284
rect 6012 18281 6040 18312
rect 6638 18300 6644 18312
rect 6696 18300 6702 18352
rect 7098 18300 7104 18352
rect 7156 18300 7162 18352
rect 5629 18275 5687 18281
rect 5629 18272 5641 18275
rect 5592 18244 5641 18272
rect 5592 18232 5598 18244
rect 5629 18241 5641 18244
rect 5675 18241 5687 18275
rect 5629 18235 5687 18241
rect 5997 18275 6055 18281
rect 5997 18241 6009 18275
rect 6043 18241 6055 18275
rect 5997 18235 6055 18241
rect 7926 18232 7932 18284
rect 7984 18272 7990 18284
rect 8665 18275 8723 18281
rect 8665 18272 8677 18275
rect 7984 18244 8677 18272
rect 7984 18232 7990 18244
rect 8665 18241 8677 18244
rect 8711 18241 8723 18275
rect 8665 18235 8723 18241
rect 8941 18275 8999 18281
rect 8941 18241 8953 18275
rect 8987 18272 8999 18275
rect 9122 18272 9128 18284
rect 8987 18244 9128 18272
rect 8987 18241 8999 18244
rect 8941 18235 8999 18241
rect 9122 18232 9128 18244
rect 9180 18232 9186 18284
rect 9950 18232 9956 18284
rect 10008 18272 10014 18284
rect 10229 18275 10287 18281
rect 10229 18272 10241 18275
rect 10008 18244 10241 18272
rect 10008 18232 10014 18244
rect 10229 18241 10241 18244
rect 10275 18241 10287 18275
rect 10229 18235 10287 18241
rect 11054 18232 11060 18284
rect 11112 18232 11118 18284
rect 11146 18232 11152 18284
rect 11204 18232 11210 18284
rect 12158 18232 12164 18284
rect 12216 18272 12222 18284
rect 12253 18275 12311 18281
rect 12253 18272 12265 18275
rect 12216 18244 12265 18272
rect 12216 18232 12222 18244
rect 12253 18241 12265 18244
rect 12299 18241 12311 18275
rect 12253 18235 12311 18241
rect 13262 18232 13268 18284
rect 13320 18272 13326 18284
rect 13541 18275 13599 18281
rect 13541 18272 13553 18275
rect 13320 18244 13553 18272
rect 13320 18232 13326 18244
rect 13541 18241 13553 18244
rect 13587 18241 13599 18275
rect 13541 18235 13599 18241
rect 14366 18232 14372 18284
rect 14424 18272 14430 18284
rect 14461 18275 14519 18281
rect 14461 18272 14473 18275
rect 14424 18244 14473 18272
rect 14424 18232 14430 18244
rect 14461 18241 14473 18244
rect 14507 18241 14519 18275
rect 14461 18235 14519 18241
rect 15470 18232 15476 18284
rect 15528 18272 15534 18284
rect 15749 18275 15807 18281
rect 15749 18272 15761 18275
rect 15528 18244 15761 18272
rect 15528 18232 15534 18244
rect 15749 18241 15761 18244
rect 15795 18241 15807 18275
rect 15749 18235 15807 18241
rect 16574 18232 16580 18284
rect 16632 18272 16638 18284
rect 16853 18275 16911 18281
rect 16853 18272 16865 18275
rect 16632 18244 16865 18272
rect 16632 18232 16638 18244
rect 16853 18241 16865 18244
rect 16899 18241 16911 18275
rect 16853 18235 16911 18241
rect 17497 18275 17555 18281
rect 17497 18241 17509 18275
rect 17543 18272 17555 18275
rect 17678 18272 17684 18284
rect 17543 18244 17684 18272
rect 17543 18241 17555 18244
rect 17497 18235 17555 18241
rect 17678 18232 17684 18244
rect 17736 18232 17742 18284
rect 3510 18204 3516 18216
rect 1872 18176 3516 18204
rect 3510 18164 3516 18176
rect 3568 18164 3574 18216
rect 6362 18164 6368 18216
rect 6420 18164 6426 18216
rect 6641 18207 6699 18213
rect 6641 18204 6653 18207
rect 6472 18176 6653 18204
rect 4709 18139 4767 18145
rect 4709 18105 4721 18139
rect 4755 18136 4767 18139
rect 6472 18136 6500 18176
rect 6641 18173 6653 18176
rect 6687 18173 6699 18207
rect 6641 18167 6699 18173
rect 8389 18207 8447 18213
rect 8389 18173 8401 18207
rect 8435 18204 8447 18207
rect 11974 18204 11980 18216
rect 8435 18176 11980 18204
rect 8435 18173 8447 18176
rect 8389 18167 8447 18173
rect 11974 18164 11980 18176
rect 12032 18164 12038 18216
rect 12158 18136 12164 18148
rect 4755 18108 6500 18136
rect 8404 18108 12164 18136
rect 4755 18105 4767 18108
rect 4709 18099 4767 18105
rect 1578 18028 1584 18080
rect 1636 18028 1642 18080
rect 3605 18071 3663 18077
rect 3605 18037 3617 18071
rect 3651 18068 3663 18071
rect 4890 18068 4896 18080
rect 3651 18040 4896 18068
rect 3651 18037 3663 18040
rect 3605 18031 3663 18037
rect 4890 18028 4896 18040
rect 4948 18028 4954 18080
rect 6181 18071 6239 18077
rect 6181 18037 6193 18071
rect 6227 18068 6239 18071
rect 8404 18068 8432 18108
rect 12158 18096 12164 18108
rect 12216 18096 12222 18148
rect 6227 18040 8432 18068
rect 6227 18037 6239 18040
rect 6181 18031 6239 18037
rect 8478 18028 8484 18080
rect 8536 18028 8542 18080
rect 9125 18071 9183 18077
rect 9125 18037 9137 18071
rect 9171 18068 9183 18071
rect 9950 18068 9956 18080
rect 9171 18040 9956 18068
rect 9171 18037 9183 18040
rect 9125 18031 9183 18037
rect 9950 18028 9956 18040
rect 10008 18028 10014 18080
rect 10042 18028 10048 18080
rect 10100 18028 10106 18080
rect 10965 18071 11023 18077
rect 10965 18037 10977 18071
rect 11011 18068 11023 18071
rect 11054 18068 11060 18080
rect 11011 18040 11060 18068
rect 11011 18037 11023 18040
rect 10965 18031 11023 18037
rect 11054 18028 11060 18040
rect 11112 18028 11118 18080
rect 11333 18071 11391 18077
rect 11333 18037 11345 18071
rect 11379 18068 11391 18071
rect 11790 18068 11796 18080
rect 11379 18040 11796 18068
rect 11379 18037 11391 18040
rect 11333 18031 11391 18037
rect 11790 18028 11796 18040
rect 11848 18028 11854 18080
rect 12434 18028 12440 18080
rect 12492 18028 12498 18080
rect 13262 18028 13268 18080
rect 13320 18068 13326 18080
rect 13357 18071 13415 18077
rect 13357 18068 13369 18071
rect 13320 18040 13369 18068
rect 13320 18028 13326 18040
rect 13357 18037 13369 18040
rect 13403 18037 13415 18071
rect 13357 18031 13415 18037
rect 14645 18071 14703 18077
rect 14645 18037 14657 18071
rect 14691 18068 14703 18071
rect 15470 18068 15476 18080
rect 14691 18040 15476 18068
rect 14691 18037 14703 18040
rect 14645 18031 14703 18037
rect 15470 18028 15476 18040
rect 15528 18028 15534 18080
rect 15562 18028 15568 18080
rect 15620 18028 15626 18080
rect 16022 18028 16028 18080
rect 16080 18068 16086 18080
rect 16669 18071 16727 18077
rect 16669 18068 16681 18071
rect 16080 18040 16681 18068
rect 16080 18028 16086 18040
rect 16669 18037 16681 18040
rect 16715 18037 16727 18071
rect 16669 18031 16727 18037
rect 17218 18028 17224 18080
rect 17276 18068 17282 18080
rect 17313 18071 17371 18077
rect 17313 18068 17325 18071
rect 17276 18040 17325 18068
rect 17276 18028 17282 18040
rect 17313 18037 17325 18040
rect 17359 18037 17371 18071
rect 17313 18031 17371 18037
rect 1104 17978 17848 18000
rect 1104 17926 1918 17978
rect 1970 17926 1982 17978
rect 2034 17926 2046 17978
rect 2098 17926 2110 17978
rect 2162 17926 2174 17978
rect 2226 17926 2238 17978
rect 2290 17926 7918 17978
rect 7970 17926 7982 17978
rect 8034 17926 8046 17978
rect 8098 17926 8110 17978
rect 8162 17926 8174 17978
rect 8226 17926 8238 17978
rect 8290 17926 13918 17978
rect 13970 17926 13982 17978
rect 14034 17926 14046 17978
rect 14098 17926 14110 17978
rect 14162 17926 14174 17978
rect 14226 17926 14238 17978
rect 14290 17926 17848 17978
rect 1104 17904 17848 17926
rect 9033 17799 9091 17805
rect 9033 17796 9045 17799
rect 8128 17768 9045 17796
rect 1397 17731 1455 17737
rect 1397 17697 1409 17731
rect 1443 17728 1455 17731
rect 4062 17728 4068 17740
rect 1443 17700 4068 17728
rect 1443 17697 1455 17700
rect 1397 17691 1455 17697
rect 4062 17688 4068 17700
rect 4120 17728 4126 17740
rect 4617 17731 4675 17737
rect 4617 17728 4629 17731
rect 4120 17700 4629 17728
rect 4120 17688 4126 17700
rect 4617 17697 4629 17700
rect 4663 17728 4675 17731
rect 6362 17728 6368 17740
rect 4663 17700 6368 17728
rect 4663 17697 4675 17700
rect 4617 17691 4675 17697
rect 6362 17688 6368 17700
rect 6420 17728 6426 17740
rect 6733 17731 6791 17737
rect 6733 17728 6745 17731
rect 6420 17700 6745 17728
rect 6420 17688 6426 17700
rect 6733 17697 6745 17700
rect 6779 17697 6791 17731
rect 6733 17691 6791 17697
rect 7006 17688 7012 17740
rect 7064 17688 7070 17740
rect 3973 17663 4031 17669
rect 3973 17660 3985 17663
rect 3804 17632 3985 17660
rect 1578 17552 1584 17604
rect 1636 17592 1642 17604
rect 1673 17595 1731 17601
rect 1673 17592 1685 17595
rect 1636 17564 1685 17592
rect 1636 17552 1642 17564
rect 1673 17561 1685 17564
rect 1719 17561 1731 17595
rect 1673 17555 1731 17561
rect 2222 17552 2228 17604
rect 2280 17552 2286 17604
rect 3234 17552 3240 17604
rect 3292 17592 3298 17604
rect 3421 17595 3479 17601
rect 3421 17592 3433 17595
rect 3292 17564 3433 17592
rect 3292 17552 3298 17564
rect 3421 17561 3433 17564
rect 3467 17561 3479 17595
rect 3421 17555 3479 17561
rect 2498 17484 2504 17536
rect 2556 17524 2562 17536
rect 3804 17524 3832 17632
rect 3973 17629 3985 17632
rect 4019 17660 4031 17663
rect 4525 17663 4583 17669
rect 4525 17660 4537 17663
rect 4019 17632 4537 17660
rect 4019 17629 4031 17632
rect 3973 17623 4031 17629
rect 4525 17629 4537 17632
rect 4571 17629 4583 17663
rect 8128 17646 8156 17768
rect 9033 17765 9045 17768
rect 9079 17765 9091 17799
rect 9033 17759 9091 17765
rect 8680 17700 9168 17728
rect 4525 17623 4583 17629
rect 2556 17496 3832 17524
rect 2556 17484 2562 17496
rect 3878 17484 3884 17536
rect 3936 17484 3942 17536
rect 4430 17484 4436 17536
rect 4488 17484 4494 17536
rect 4540 17524 4568 17623
rect 4890 17552 4896 17604
rect 4948 17552 4954 17604
rect 6454 17592 6460 17604
rect 6118 17564 6460 17592
rect 6454 17552 6460 17564
rect 6512 17552 6518 17604
rect 6638 17552 6644 17604
rect 6696 17552 6702 17604
rect 6546 17524 6552 17536
rect 4540 17496 6552 17524
rect 6546 17484 6552 17496
rect 6604 17524 6610 17536
rect 8680 17524 8708 17700
rect 9140 17672 9168 17700
rect 9766 17688 9772 17740
rect 9824 17688 9830 17740
rect 10042 17688 10048 17740
rect 10100 17688 10106 17740
rect 11885 17731 11943 17737
rect 11885 17697 11897 17731
rect 11931 17728 11943 17731
rect 13538 17728 13544 17740
rect 11931 17700 13544 17728
rect 11931 17697 11943 17700
rect 11885 17691 11943 17697
rect 13538 17688 13544 17700
rect 13596 17728 13602 17740
rect 14645 17731 14703 17737
rect 14645 17728 14657 17731
rect 13596 17700 14657 17728
rect 13596 17688 13602 17700
rect 14645 17697 14657 17700
rect 14691 17697 14703 17731
rect 14645 17691 14703 17697
rect 14921 17731 14979 17737
rect 14921 17697 14933 17731
rect 14967 17728 14979 17731
rect 15562 17728 15568 17740
rect 14967 17700 15568 17728
rect 14967 17697 14979 17700
rect 14921 17691 14979 17697
rect 15562 17688 15568 17700
rect 15620 17688 15626 17740
rect 9122 17620 9128 17672
rect 9180 17620 9186 17672
rect 14277 17663 14335 17669
rect 14277 17660 14289 17663
rect 14108 17632 14289 17660
rect 8757 17595 8815 17601
rect 8757 17561 8769 17595
rect 8803 17561 8815 17595
rect 8757 17555 8815 17561
rect 6604 17496 8708 17524
rect 8772 17524 8800 17555
rect 11054 17552 11060 17604
rect 11112 17552 11118 17604
rect 11422 17552 11428 17604
rect 11480 17592 11486 17604
rect 11793 17595 11851 17601
rect 11793 17592 11805 17595
rect 11480 17564 11805 17592
rect 11480 17552 11486 17564
rect 11793 17561 11805 17564
rect 11839 17561 11851 17595
rect 11793 17555 11851 17561
rect 12158 17552 12164 17604
rect 12216 17552 12222 17604
rect 12618 17552 12624 17604
rect 12676 17552 12682 17604
rect 13446 17552 13452 17604
rect 13504 17592 13510 17604
rect 13909 17595 13967 17601
rect 13909 17592 13921 17595
rect 13504 17564 13921 17592
rect 13504 17552 13510 17564
rect 13909 17561 13921 17564
rect 13955 17561 13967 17595
rect 13909 17555 13967 17561
rect 12250 17524 12256 17536
rect 8772 17496 12256 17524
rect 6604 17484 6610 17496
rect 12250 17484 12256 17496
rect 12308 17484 12314 17536
rect 12342 17484 12348 17536
rect 12400 17524 12406 17536
rect 14108 17524 14136 17632
rect 14277 17629 14289 17632
rect 14323 17660 14335 17663
rect 14550 17660 14556 17672
rect 14323 17632 14556 17660
rect 14323 17629 14335 17632
rect 14277 17623 14335 17629
rect 14550 17620 14556 17632
rect 14608 17620 14614 17672
rect 16758 17620 16764 17672
rect 16816 17660 16822 17672
rect 16853 17663 16911 17669
rect 16853 17660 16865 17663
rect 16816 17632 16865 17660
rect 16816 17620 16822 17632
rect 16853 17629 16865 17632
rect 16899 17629 16911 17663
rect 16853 17623 16911 17629
rect 15654 17552 15660 17604
rect 15712 17552 15718 17604
rect 16482 17552 16488 17604
rect 16540 17592 16546 17604
rect 16669 17595 16727 17601
rect 16669 17592 16681 17595
rect 16540 17564 16681 17592
rect 16540 17552 16546 17564
rect 16669 17561 16681 17564
rect 16715 17561 16727 17595
rect 16669 17555 16727 17561
rect 12400 17496 14136 17524
rect 14185 17527 14243 17533
rect 12400 17484 12406 17496
rect 14185 17493 14197 17527
rect 14231 17524 14243 17527
rect 14274 17524 14280 17536
rect 14231 17496 14280 17524
rect 14231 17493 14243 17496
rect 14185 17487 14243 17493
rect 14274 17484 14280 17496
rect 14332 17484 14338 17536
rect 16945 17527 17003 17533
rect 16945 17493 16957 17527
rect 16991 17524 17003 17527
rect 17034 17524 17040 17536
rect 16991 17496 17040 17524
rect 16991 17493 17003 17496
rect 16945 17487 17003 17493
rect 17034 17484 17040 17496
rect 17092 17484 17098 17536
rect 1104 17434 17848 17456
rect 1104 17382 2658 17434
rect 2710 17382 2722 17434
rect 2774 17382 2786 17434
rect 2838 17382 2850 17434
rect 2902 17382 2914 17434
rect 2966 17382 2978 17434
rect 3030 17382 8658 17434
rect 8710 17382 8722 17434
rect 8774 17382 8786 17434
rect 8838 17382 8850 17434
rect 8902 17382 8914 17434
rect 8966 17382 8978 17434
rect 9030 17382 14658 17434
rect 14710 17382 14722 17434
rect 14774 17382 14786 17434
rect 14838 17382 14850 17434
rect 14902 17382 14914 17434
rect 14966 17382 14978 17434
rect 15030 17382 17848 17434
rect 1104 17360 17848 17382
rect 1302 17280 1308 17332
rect 1360 17320 1366 17332
rect 1397 17323 1455 17329
rect 1397 17320 1409 17323
rect 1360 17292 1409 17320
rect 1360 17280 1366 17292
rect 1397 17289 1409 17292
rect 1443 17289 1455 17323
rect 1397 17283 1455 17289
rect 2222 17280 2228 17332
rect 2280 17280 2286 17332
rect 3510 17280 3516 17332
rect 3568 17280 3574 17332
rect 6454 17280 6460 17332
rect 6512 17280 6518 17332
rect 7098 17280 7104 17332
rect 7156 17280 7162 17332
rect 9122 17280 9128 17332
rect 9180 17320 9186 17332
rect 11146 17320 11152 17332
rect 9180 17292 11152 17320
rect 9180 17280 9186 17292
rect 4430 17212 4436 17264
rect 4488 17212 4494 17264
rect 8205 17255 8263 17261
rect 8205 17221 8217 17255
rect 8251 17252 8263 17255
rect 8478 17252 8484 17264
rect 8251 17224 8484 17252
rect 8251 17221 8263 17224
rect 8205 17215 8263 17221
rect 8478 17212 8484 17224
rect 8536 17212 8542 17264
rect 9214 17212 9220 17264
rect 9272 17212 9278 17264
rect 1581 17187 1639 17193
rect 1581 17153 1593 17187
rect 1627 17153 1639 17187
rect 1581 17147 1639 17153
rect 2133 17187 2191 17193
rect 2133 17153 2145 17187
rect 2179 17184 2191 17187
rect 2498 17184 2504 17196
rect 2179 17156 2504 17184
rect 2179 17153 2191 17156
rect 2133 17147 2191 17153
rect 1596 17116 1624 17147
rect 2498 17144 2504 17156
rect 2556 17144 2562 17196
rect 6546 17144 6552 17196
rect 6604 17184 6610 17196
rect 10888 17193 10916 17292
rect 11146 17280 11152 17292
rect 11204 17280 11210 17332
rect 12529 17323 12587 17329
rect 12529 17289 12541 17323
rect 12575 17320 12587 17323
rect 12618 17320 12624 17332
rect 12575 17292 12624 17320
rect 12575 17289 12587 17292
rect 12529 17283 12587 17289
rect 12618 17280 12624 17292
rect 12676 17280 12682 17332
rect 15654 17280 15660 17332
rect 15712 17280 15718 17332
rect 13538 17252 13544 17264
rect 13004 17224 13544 17252
rect 7009 17187 7067 17193
rect 7009 17184 7021 17187
rect 6604 17156 7021 17184
rect 6604 17144 6610 17156
rect 7009 17153 7021 17156
rect 7055 17153 7067 17187
rect 7009 17147 7067 17153
rect 10873 17187 10931 17193
rect 10873 17153 10885 17187
rect 10919 17184 10931 17187
rect 12342 17184 12348 17196
rect 10919 17156 12348 17184
rect 10919 17153 10931 17156
rect 10873 17147 10931 17153
rect 12342 17144 12348 17156
rect 12400 17184 12406 17196
rect 13004 17193 13032 17224
rect 13538 17212 13544 17224
rect 13596 17212 13602 17264
rect 14274 17212 14280 17264
rect 14332 17212 14338 17264
rect 12437 17187 12495 17193
rect 12437 17184 12449 17187
rect 12400 17156 12449 17184
rect 12400 17144 12406 17156
rect 12437 17153 12449 17156
rect 12483 17153 12495 17187
rect 12437 17147 12495 17153
rect 12989 17187 13047 17193
rect 12989 17153 13001 17187
rect 13035 17153 13047 17187
rect 12989 17147 13047 17153
rect 14550 17144 14556 17196
rect 14608 17184 14614 17196
rect 15565 17187 15623 17193
rect 15565 17184 15577 17187
rect 14608 17156 15577 17184
rect 14608 17144 14614 17156
rect 15565 17153 15577 17156
rect 15611 17184 15623 17187
rect 16758 17184 16764 17196
rect 15611 17156 16764 17184
rect 15611 17153 15623 17156
rect 15565 17147 15623 17153
rect 16758 17144 16764 17156
rect 16816 17144 16822 17196
rect 3050 17116 3056 17128
rect 1596 17088 3056 17116
rect 3050 17076 3056 17088
rect 3108 17076 3114 17128
rect 4246 17076 4252 17128
rect 4304 17116 4310 17128
rect 4985 17119 5043 17125
rect 4985 17116 4997 17119
rect 4304 17088 4997 17116
rect 4304 17076 4310 17088
rect 4985 17085 4997 17088
rect 5031 17085 5043 17119
rect 4985 17079 5043 17085
rect 5261 17119 5319 17125
rect 5261 17085 5273 17119
rect 5307 17085 5319 17119
rect 5261 17079 5319 17085
rect 7929 17119 7987 17125
rect 7929 17085 7941 17119
rect 7975 17116 7987 17119
rect 9858 17116 9864 17128
rect 7975 17088 9864 17116
rect 7975 17085 7987 17088
rect 7929 17079 7987 17085
rect 3970 16940 3976 16992
rect 4028 16980 4034 16992
rect 5276 16980 5304 17079
rect 9858 17076 9864 17088
rect 9916 17076 9922 17128
rect 9953 17119 10011 17125
rect 9953 17085 9965 17119
rect 9999 17116 10011 17119
rect 12066 17116 12072 17128
rect 9999 17088 12072 17116
rect 9999 17085 10011 17088
rect 9953 17079 10011 17085
rect 12066 17076 12072 17088
rect 12124 17076 12130 17128
rect 13262 17076 13268 17128
rect 13320 17076 13326 17128
rect 15013 17119 15071 17125
rect 15013 17085 15025 17119
rect 15059 17116 15071 17119
rect 16850 17116 16856 17128
rect 15059 17088 16856 17116
rect 15059 17085 15071 17088
rect 15013 17079 15071 17085
rect 16850 17076 16856 17088
rect 16908 17076 16914 17128
rect 4028 16952 5304 16980
rect 10965 16983 11023 16989
rect 4028 16940 4034 16952
rect 10965 16949 10977 16983
rect 11011 16980 11023 16983
rect 11146 16980 11152 16992
rect 11011 16952 11152 16980
rect 11011 16949 11023 16952
rect 10965 16943 11023 16949
rect 11146 16940 11152 16952
rect 11204 16940 11210 16992
rect 1104 16890 17848 16912
rect 1104 16838 1918 16890
rect 1970 16838 1982 16890
rect 2034 16838 2046 16890
rect 2098 16838 2110 16890
rect 2162 16838 2174 16890
rect 2226 16838 2238 16890
rect 2290 16838 7918 16890
rect 7970 16838 7982 16890
rect 8034 16838 8046 16890
rect 8098 16838 8110 16890
rect 8162 16838 8174 16890
rect 8226 16838 8238 16890
rect 8290 16838 13918 16890
rect 13970 16838 13982 16890
rect 14034 16838 14046 16890
rect 14098 16838 14110 16890
rect 14162 16838 14174 16890
rect 14226 16838 14238 16890
rect 14290 16838 17848 16890
rect 1104 16816 17848 16838
rect 3421 16779 3479 16785
rect 3421 16745 3433 16779
rect 3467 16776 3479 16779
rect 4338 16776 4344 16788
rect 3467 16748 4344 16776
rect 3467 16745 3479 16748
rect 3421 16739 3479 16745
rect 4338 16736 4344 16748
rect 4396 16736 4402 16788
rect 9125 16779 9183 16785
rect 9125 16745 9137 16779
rect 9171 16776 9183 16779
rect 9214 16776 9220 16788
rect 9171 16748 9220 16776
rect 9171 16745 9183 16748
rect 9125 16739 9183 16745
rect 9214 16736 9220 16748
rect 9272 16736 9278 16788
rect 9950 16736 9956 16788
rect 10008 16776 10014 16788
rect 10118 16779 10176 16785
rect 10118 16776 10130 16779
rect 10008 16748 10130 16776
rect 10008 16736 10014 16748
rect 10118 16745 10130 16748
rect 10164 16745 10176 16779
rect 10118 16739 10176 16745
rect 3344 16680 4200 16708
rect 3344 16652 3372 16680
rect 3145 16643 3203 16649
rect 3145 16609 3157 16643
rect 3191 16640 3203 16643
rect 3326 16640 3332 16652
rect 3191 16612 3332 16640
rect 3191 16609 3203 16612
rect 3145 16603 3203 16609
rect 3326 16600 3332 16612
rect 3384 16600 3390 16652
rect 1394 16532 1400 16584
rect 1452 16572 1458 16584
rect 1581 16575 1639 16581
rect 1581 16572 1593 16575
rect 1452 16544 1593 16572
rect 1452 16532 1458 16544
rect 1581 16541 1593 16544
rect 1627 16541 1639 16575
rect 1581 16535 1639 16541
rect 3053 16575 3111 16581
rect 3053 16541 3065 16575
rect 3099 16572 3111 16575
rect 4062 16572 4068 16584
rect 3099 16544 4068 16572
rect 3099 16541 3111 16544
rect 3053 16535 3111 16541
rect 4062 16532 4068 16544
rect 4120 16532 4126 16584
rect 4172 16581 4200 16680
rect 13906 16668 13912 16720
rect 13964 16708 13970 16720
rect 15197 16711 15255 16717
rect 15197 16708 15209 16711
rect 13964 16680 15209 16708
rect 13964 16668 13970 16680
rect 15197 16677 15209 16680
rect 15243 16677 15255 16711
rect 15197 16671 15255 16677
rect 5810 16640 5816 16652
rect 4448 16612 5816 16640
rect 4448 16581 4476 16612
rect 5810 16600 5816 16612
rect 5868 16600 5874 16652
rect 9122 16600 9128 16652
rect 9180 16640 9186 16652
rect 9180 16612 9260 16640
rect 9180 16600 9186 16612
rect 9232 16581 9260 16612
rect 9858 16600 9864 16652
rect 9916 16640 9922 16652
rect 10134 16640 10140 16652
rect 9916 16612 10140 16640
rect 9916 16600 9922 16612
rect 10134 16600 10140 16612
rect 10192 16600 10198 16652
rect 13538 16600 13544 16652
rect 13596 16640 13602 16652
rect 15749 16643 15807 16649
rect 15749 16640 15761 16643
rect 13596 16612 15761 16640
rect 13596 16600 13602 16612
rect 15749 16609 15761 16612
rect 15795 16609 15807 16643
rect 15749 16603 15807 16609
rect 16022 16600 16028 16652
rect 16080 16600 16086 16652
rect 4157 16575 4215 16581
rect 4157 16541 4169 16575
rect 4203 16541 4215 16575
rect 4157 16535 4215 16541
rect 4249 16575 4307 16581
rect 4249 16541 4261 16575
rect 4295 16541 4307 16575
rect 4249 16535 4307 16541
rect 4433 16575 4491 16581
rect 4433 16541 4445 16575
rect 4479 16541 4491 16575
rect 4433 16535 4491 16541
rect 9217 16575 9275 16581
rect 9217 16541 9229 16575
rect 9263 16541 9275 16575
rect 9217 16535 9275 16541
rect 842 16396 848 16448
rect 900 16436 906 16448
rect 1397 16439 1455 16445
rect 1397 16436 1409 16439
rect 900 16408 1409 16436
rect 900 16396 906 16408
rect 1397 16405 1409 16408
rect 1443 16405 1455 16439
rect 1397 16399 1455 16405
rect 3789 16439 3847 16445
rect 3789 16405 3801 16439
rect 3835 16436 3847 16439
rect 4154 16436 4160 16448
rect 3835 16408 4160 16436
rect 3835 16405 3847 16408
rect 3789 16399 3847 16405
rect 4154 16396 4160 16408
rect 4212 16396 4218 16448
rect 4264 16436 4292 16535
rect 12986 16532 12992 16584
rect 13044 16532 13050 16584
rect 13265 16575 13323 16581
rect 13265 16541 13277 16575
rect 13311 16572 13323 16575
rect 13906 16572 13912 16584
rect 13311 16544 13912 16572
rect 13311 16541 13323 16544
rect 13265 16535 13323 16541
rect 13906 16532 13912 16544
rect 13964 16532 13970 16584
rect 14921 16575 14979 16581
rect 14921 16541 14933 16575
rect 14967 16541 14979 16575
rect 14921 16535 14979 16541
rect 15105 16575 15163 16581
rect 15105 16541 15117 16575
rect 15151 16572 15163 16575
rect 15381 16575 15439 16581
rect 15381 16572 15393 16575
rect 15151 16544 15393 16572
rect 15151 16541 15163 16544
rect 15105 16535 15163 16541
rect 15381 16541 15393 16544
rect 15427 16541 15439 16575
rect 15381 16535 15439 16541
rect 11146 16464 11152 16516
rect 11204 16464 11210 16516
rect 11885 16507 11943 16513
rect 11885 16473 11897 16507
rect 11931 16504 11943 16507
rect 12434 16504 12440 16516
rect 11931 16476 12440 16504
rect 11931 16473 11943 16476
rect 11885 16467 11943 16473
rect 12434 16464 12440 16476
rect 12492 16464 12498 16516
rect 14936 16504 14964 16535
rect 15396 16504 15424 16535
rect 15562 16532 15568 16584
rect 15620 16532 15626 16584
rect 14936 16476 15332 16504
rect 15396 16476 15884 16504
rect 6546 16436 6552 16448
rect 4264 16408 6552 16436
rect 6546 16396 6552 16408
rect 6604 16396 6610 16448
rect 12802 16396 12808 16448
rect 12860 16396 12866 16448
rect 13173 16439 13231 16445
rect 13173 16405 13185 16439
rect 13219 16436 13231 16439
rect 13446 16436 13452 16448
rect 13219 16408 13452 16436
rect 13219 16405 13231 16408
rect 13173 16399 13231 16405
rect 13446 16396 13452 16408
rect 13504 16396 13510 16448
rect 15013 16439 15071 16445
rect 15013 16405 15025 16439
rect 15059 16436 15071 16439
rect 15102 16436 15108 16448
rect 15059 16408 15108 16436
rect 15059 16405 15071 16408
rect 15013 16399 15071 16405
rect 15102 16396 15108 16408
rect 15160 16396 15166 16448
rect 15304 16436 15332 16476
rect 15856 16448 15884 16476
rect 17034 16464 17040 16516
rect 17092 16464 17098 16516
rect 15562 16436 15568 16448
rect 15304 16408 15568 16436
rect 15562 16396 15568 16408
rect 15620 16396 15626 16448
rect 15838 16396 15844 16448
rect 15896 16436 15902 16448
rect 17497 16439 17555 16445
rect 17497 16436 17509 16439
rect 15896 16408 17509 16436
rect 15896 16396 15902 16408
rect 17497 16405 17509 16408
rect 17543 16405 17555 16439
rect 17497 16399 17555 16405
rect 1104 16346 17848 16368
rect 1104 16294 2658 16346
rect 2710 16294 2722 16346
rect 2774 16294 2786 16346
rect 2838 16294 2850 16346
rect 2902 16294 2914 16346
rect 2966 16294 2978 16346
rect 3030 16294 8658 16346
rect 8710 16294 8722 16346
rect 8774 16294 8786 16346
rect 8838 16294 8850 16346
rect 8902 16294 8914 16346
rect 8966 16294 8978 16346
rect 9030 16294 14658 16346
rect 14710 16294 14722 16346
rect 14774 16294 14786 16346
rect 14838 16294 14850 16346
rect 14902 16294 14914 16346
rect 14966 16294 14978 16346
rect 15030 16294 17848 16346
rect 1104 16272 17848 16294
rect 2869 16235 2927 16241
rect 2869 16201 2881 16235
rect 2915 16232 2927 16235
rect 3050 16232 3056 16244
rect 2915 16204 3056 16232
rect 2915 16201 2927 16204
rect 2869 16195 2927 16201
rect 3050 16192 3056 16204
rect 3108 16192 3114 16244
rect 4062 16192 4068 16244
rect 4120 16232 4126 16244
rect 5169 16235 5227 16241
rect 5169 16232 5181 16235
rect 4120 16204 5181 16232
rect 4120 16192 4126 16204
rect 5169 16201 5181 16204
rect 5215 16201 5227 16235
rect 5169 16195 5227 16201
rect 5810 16192 5816 16244
rect 5868 16192 5874 16244
rect 7282 16192 7288 16244
rect 7340 16232 7346 16244
rect 7834 16232 7840 16244
rect 7340 16204 7840 16232
rect 7340 16192 7346 16204
rect 7834 16192 7840 16204
rect 7892 16232 7898 16244
rect 8757 16235 8815 16241
rect 8757 16232 8769 16235
rect 7892 16204 8769 16232
rect 7892 16192 7898 16204
rect 8757 16201 8769 16204
rect 8803 16201 8815 16235
rect 8757 16195 8815 16201
rect 12342 16192 12348 16244
rect 12400 16232 12406 16244
rect 13998 16232 14004 16244
rect 12400 16204 14004 16232
rect 12400 16192 12406 16204
rect 3878 16124 3884 16176
rect 3936 16124 3942 16176
rect 4338 16124 4344 16176
rect 4396 16124 4402 16176
rect 7377 16167 7435 16173
rect 7377 16164 7389 16167
rect 5828 16136 6500 16164
rect 1578 16056 1584 16108
rect 1636 16056 1642 16108
rect 2133 16099 2191 16105
rect 2133 16065 2145 16099
rect 2179 16096 2191 16099
rect 2498 16096 2504 16108
rect 2179 16068 2504 16096
rect 2179 16065 2191 16068
rect 2133 16059 2191 16065
rect 2498 16056 2504 16068
rect 2556 16056 2562 16108
rect 5828 16105 5856 16136
rect 5537 16099 5595 16105
rect 5537 16065 5549 16099
rect 5583 16096 5595 16099
rect 5813 16099 5871 16105
rect 5813 16096 5825 16099
rect 5583 16068 5825 16096
rect 5583 16065 5595 16068
rect 5537 16059 5595 16065
rect 5813 16065 5825 16068
rect 5859 16065 5871 16099
rect 5813 16059 5871 16065
rect 5997 16099 6055 16105
rect 5997 16065 6009 16099
rect 6043 16096 6055 16099
rect 6365 16099 6423 16105
rect 6365 16096 6377 16099
rect 6043 16068 6377 16096
rect 6043 16065 6055 16068
rect 5997 16059 6055 16065
rect 6365 16065 6377 16068
rect 6411 16065 6423 16099
rect 6365 16059 6423 16065
rect 3142 15988 3148 16040
rect 3200 16028 3206 16040
rect 3970 16028 3976 16040
rect 3200 16000 3976 16028
rect 3200 15988 3206 16000
rect 3970 15988 3976 16000
rect 4028 16028 4034 16040
rect 4617 16031 4675 16037
rect 4617 16028 4629 16031
rect 4028 16000 4629 16028
rect 4028 15988 4034 16000
rect 4617 15997 4629 16000
rect 4663 15997 4675 16031
rect 4617 15991 4675 15997
rect 5629 16031 5687 16037
rect 5629 15997 5641 16031
rect 5675 16028 5687 16031
rect 6012 16028 6040 16059
rect 5675 16000 6040 16028
rect 5675 15997 5687 16000
rect 5629 15991 5687 15997
rect 6472 15960 6500 16136
rect 6564 16136 7389 16164
rect 6564 16108 6592 16136
rect 7377 16133 7389 16136
rect 7423 16133 7435 16167
rect 9582 16164 9588 16176
rect 7377 16127 7435 16133
rect 8680 16136 9588 16164
rect 6546 16056 6552 16108
rect 6604 16056 6610 16108
rect 7009 16099 7067 16105
rect 7009 16065 7021 16099
rect 7055 16096 7067 16099
rect 7098 16096 7104 16108
rect 7055 16068 7104 16096
rect 7055 16065 7067 16068
rect 7009 16059 7067 16065
rect 7098 16056 7104 16068
rect 7156 16056 7162 16108
rect 7193 16099 7251 16105
rect 7193 16065 7205 16099
rect 7239 16065 7251 16099
rect 7193 16059 7251 16065
rect 6733 16031 6791 16037
rect 6733 15997 6745 16031
rect 6779 16028 6791 16031
rect 6825 16031 6883 16037
rect 6825 16028 6837 16031
rect 6779 16000 6837 16028
rect 6779 15997 6791 16000
rect 6733 15991 6791 15997
rect 6825 15997 6837 16000
rect 6871 15997 6883 16031
rect 7208 16028 7236 16059
rect 7282 16056 7288 16108
rect 7340 16056 7346 16108
rect 8680 16105 8708 16136
rect 9582 16124 9588 16136
rect 9640 16124 9646 16176
rect 12526 16164 12532 16176
rect 12452 16136 12532 16164
rect 7469 16099 7527 16105
rect 7469 16065 7481 16099
rect 7515 16065 7527 16099
rect 7469 16059 7527 16065
rect 8665 16099 8723 16105
rect 8665 16065 8677 16099
rect 8711 16065 8723 16099
rect 8665 16059 8723 16065
rect 7484 16028 7512 16059
rect 8846 16056 8852 16108
rect 8904 16056 8910 16108
rect 12250 16056 12256 16108
rect 12308 16056 12314 16108
rect 12452 16105 12480 16136
rect 12526 16124 12532 16136
rect 12584 16124 12590 16176
rect 12636 16105 12664 16204
rect 13998 16192 14004 16204
rect 14056 16232 14062 16244
rect 14458 16232 14464 16244
rect 14056 16204 14464 16232
rect 14056 16192 14062 16204
rect 14458 16192 14464 16204
rect 14516 16192 14522 16244
rect 14826 16192 14832 16244
rect 14884 16232 14890 16244
rect 15102 16232 15108 16244
rect 14884 16204 15108 16232
rect 14884 16192 14890 16204
rect 15102 16192 15108 16204
rect 15160 16192 15166 16244
rect 13357 16167 13415 16173
rect 13357 16133 13369 16167
rect 13403 16164 13415 16167
rect 14369 16167 14427 16173
rect 14369 16164 14381 16167
rect 13403 16136 14381 16164
rect 13403 16133 13415 16136
rect 13357 16127 13415 16133
rect 14369 16133 14381 16136
rect 14415 16164 14427 16167
rect 15013 16167 15071 16173
rect 15013 16164 15025 16167
rect 14415 16136 15025 16164
rect 14415 16133 14427 16136
rect 14369 16127 14427 16133
rect 15013 16133 15025 16136
rect 15059 16133 15071 16167
rect 15013 16127 15071 16133
rect 15562 16124 15568 16176
rect 15620 16164 15626 16176
rect 16482 16164 16488 16176
rect 15620 16136 16488 16164
rect 15620 16124 15626 16136
rect 12437 16099 12495 16105
rect 12437 16065 12449 16099
rect 12483 16065 12495 16099
rect 12437 16059 12495 16065
rect 12621 16099 12679 16105
rect 12621 16065 12633 16099
rect 12667 16065 12679 16099
rect 12621 16059 12679 16065
rect 12802 16056 12808 16108
rect 12860 16056 12866 16108
rect 12986 16056 12992 16108
rect 13044 16096 13050 16108
rect 13265 16099 13323 16105
rect 13265 16096 13277 16099
rect 13044 16068 13277 16096
rect 13044 16056 13050 16068
rect 13265 16065 13277 16068
rect 13311 16096 13323 16099
rect 13725 16099 13783 16105
rect 13725 16096 13737 16099
rect 13311 16068 13737 16096
rect 13311 16065 13323 16068
rect 13265 16059 13323 16065
rect 13725 16065 13737 16068
rect 13771 16065 13783 16099
rect 13725 16059 13783 16065
rect 12529 16031 12587 16037
rect 7208 16000 12434 16028
rect 6825 15991 6883 15997
rect 7742 15960 7748 15972
rect 6472 15932 7748 15960
rect 7742 15920 7748 15932
rect 7800 15920 7806 15972
rect 12406 15960 12434 16000
rect 12529 15997 12541 16031
rect 12575 16028 12587 16031
rect 13078 16028 13084 16040
rect 12575 16000 13084 16028
rect 12575 15997 12587 16000
rect 12529 15991 12587 15997
rect 13078 15988 13084 16000
rect 13136 16028 13142 16040
rect 13354 16028 13360 16040
rect 13136 16000 13360 16028
rect 13136 15988 13142 16000
rect 13354 15988 13360 16000
rect 13412 15988 13418 16040
rect 13541 16031 13599 16037
rect 13541 15997 13553 16031
rect 13587 15997 13599 16031
rect 13740 16028 13768 16059
rect 13906 16056 13912 16108
rect 13964 16056 13970 16108
rect 13998 16056 14004 16108
rect 14056 16056 14062 16108
rect 14185 16099 14243 16105
rect 14185 16065 14197 16099
rect 14231 16096 14243 16099
rect 14645 16099 14703 16105
rect 14231 16068 14596 16096
rect 14231 16065 14243 16068
rect 14185 16059 14243 16065
rect 14461 16031 14519 16037
rect 14461 16028 14473 16031
rect 13740 16000 14473 16028
rect 13541 15991 13599 15997
rect 14461 15997 14473 16000
rect 14507 15997 14519 16031
rect 14461 15991 14519 15997
rect 12897 15963 12955 15969
rect 12897 15960 12909 15963
rect 12406 15932 12909 15960
rect 12897 15929 12909 15932
rect 12943 15929 12955 15963
rect 13556 15960 13584 15991
rect 13814 15960 13820 15972
rect 13556 15932 13820 15960
rect 12897 15923 12955 15929
rect 13814 15920 13820 15932
rect 13872 15920 13878 15972
rect 14568 15960 14596 16068
rect 14645 16065 14657 16099
rect 14691 16065 14703 16099
rect 14645 16059 14703 16065
rect 14660 16028 14688 16059
rect 14826 16056 14832 16108
rect 14884 16056 14890 16108
rect 14918 16056 14924 16108
rect 14976 16056 14982 16108
rect 15672 16105 15700 16136
rect 16482 16124 16488 16136
rect 16540 16124 16546 16176
rect 15105 16099 15163 16105
rect 15105 16065 15117 16099
rect 15151 16065 15163 16099
rect 15105 16059 15163 16065
rect 15657 16099 15715 16105
rect 15657 16065 15669 16099
rect 15703 16065 15715 16099
rect 15657 16059 15715 16065
rect 14936 16028 14964 16056
rect 14660 16000 14964 16028
rect 15010 15988 15016 16040
rect 15068 16028 15074 16040
rect 15120 16028 15148 16059
rect 15838 16056 15844 16108
rect 15896 16056 15902 16108
rect 16758 16056 16764 16108
rect 16816 16096 16822 16108
rect 16853 16099 16911 16105
rect 16853 16096 16865 16099
rect 16816 16068 16865 16096
rect 16816 16056 16822 16068
rect 16853 16065 16865 16068
rect 16899 16065 16911 16099
rect 16853 16059 16911 16065
rect 15286 16028 15292 16040
rect 15068 16000 15292 16028
rect 15068 15988 15074 16000
rect 15286 15988 15292 16000
rect 15344 16028 15350 16040
rect 15749 16031 15807 16037
rect 15749 16028 15761 16031
rect 15344 16000 15761 16028
rect 15344 15988 15350 16000
rect 15749 15997 15761 16000
rect 15795 15997 15807 16031
rect 15749 15991 15807 15997
rect 14826 15960 14832 15972
rect 14568 15932 14832 15960
rect 14826 15920 14832 15932
rect 14884 15920 14890 15972
rect 842 15852 848 15904
rect 900 15892 906 15904
rect 1397 15895 1455 15901
rect 1397 15892 1409 15895
rect 900 15864 1409 15892
rect 900 15852 906 15864
rect 1397 15861 1409 15864
rect 1443 15861 1455 15895
rect 1397 15855 1455 15861
rect 2225 15895 2283 15901
rect 2225 15861 2237 15895
rect 2271 15892 2283 15895
rect 2314 15892 2320 15904
rect 2271 15864 2320 15892
rect 2271 15861 2283 15864
rect 2225 15855 2283 15861
rect 2314 15852 2320 15864
rect 2372 15852 2378 15904
rect 9582 15852 9588 15904
rect 9640 15892 9646 15904
rect 11698 15892 11704 15904
rect 9640 15864 11704 15892
rect 9640 15852 9646 15864
rect 11698 15852 11704 15864
rect 11756 15852 11762 15904
rect 12069 15895 12127 15901
rect 12069 15861 12081 15895
rect 12115 15892 12127 15895
rect 12158 15892 12164 15904
rect 12115 15864 12164 15892
rect 12115 15861 12127 15864
rect 12069 15855 12127 15861
rect 12158 15852 12164 15864
rect 12216 15852 12222 15904
rect 13354 15852 13360 15904
rect 13412 15892 13418 15904
rect 13725 15895 13783 15901
rect 13725 15892 13737 15895
rect 13412 15864 13737 15892
rect 13412 15852 13418 15864
rect 13725 15861 13737 15864
rect 13771 15861 13783 15895
rect 13725 15855 13783 15861
rect 16942 15852 16948 15904
rect 17000 15852 17006 15904
rect 1104 15802 17848 15824
rect 1104 15750 1918 15802
rect 1970 15750 1982 15802
rect 2034 15750 2046 15802
rect 2098 15750 2110 15802
rect 2162 15750 2174 15802
rect 2226 15750 2238 15802
rect 2290 15750 7918 15802
rect 7970 15750 7982 15802
rect 8034 15750 8046 15802
rect 8098 15750 8110 15802
rect 8162 15750 8174 15802
rect 8226 15750 8238 15802
rect 8290 15750 13918 15802
rect 13970 15750 13982 15802
rect 14034 15750 14046 15802
rect 14098 15750 14110 15802
rect 14162 15750 14174 15802
rect 14226 15750 14238 15802
rect 14290 15750 17848 15802
rect 1104 15728 17848 15750
rect 1394 15648 1400 15700
rect 1452 15648 1458 15700
rect 3326 15648 3332 15700
rect 3384 15648 3390 15700
rect 6641 15691 6699 15697
rect 6641 15688 6653 15691
rect 3620 15660 6653 15688
rect 3620 15620 3648 15660
rect 3528 15592 3648 15620
rect 3142 15444 3148 15496
rect 3200 15444 3206 15496
rect 3528 15493 3556 15592
rect 4246 15552 4252 15564
rect 3896 15524 4252 15552
rect 3513 15487 3571 15493
rect 3513 15453 3525 15487
rect 3559 15453 3571 15487
rect 3513 15447 3571 15453
rect 3605 15487 3663 15493
rect 3605 15453 3617 15487
rect 3651 15484 3663 15487
rect 3896 15484 3924 15524
rect 4246 15512 4252 15524
rect 4304 15512 4310 15564
rect 4724 15493 4752 15660
rect 6641 15657 6653 15660
rect 6687 15657 6699 15691
rect 6641 15651 6699 15657
rect 8846 15648 8852 15700
rect 8904 15688 8910 15700
rect 9493 15691 9551 15697
rect 9493 15688 9505 15691
rect 8904 15660 9505 15688
rect 8904 15648 8910 15660
rect 9493 15657 9505 15660
rect 9539 15688 9551 15691
rect 11517 15691 11575 15697
rect 11517 15688 11529 15691
rect 9539 15660 11529 15688
rect 9539 15657 9551 15660
rect 9493 15651 9551 15657
rect 11517 15657 11529 15660
rect 11563 15657 11575 15691
rect 11517 15651 11575 15657
rect 11698 15648 11704 15700
rect 11756 15688 11762 15700
rect 13541 15691 13599 15697
rect 13541 15688 13553 15691
rect 11756 15660 13553 15688
rect 11756 15648 11762 15660
rect 13541 15657 13553 15660
rect 13587 15657 13599 15691
rect 13541 15651 13599 15657
rect 13630 15648 13636 15700
rect 13688 15688 13694 15700
rect 15013 15691 15071 15697
rect 15013 15688 15025 15691
rect 13688 15660 15025 15688
rect 13688 15648 13694 15660
rect 15013 15657 15025 15660
rect 15059 15657 15071 15691
rect 15013 15651 15071 15657
rect 7006 15620 7012 15632
rect 6288 15592 7012 15620
rect 3651 15456 3924 15484
rect 4157 15487 4215 15493
rect 3651 15453 3663 15456
rect 3605 15447 3663 15453
rect 4157 15453 4169 15487
rect 4203 15484 4215 15487
rect 4433 15487 4491 15493
rect 4433 15484 4445 15487
rect 4203 15456 4445 15484
rect 4203 15453 4215 15456
rect 4157 15447 4215 15453
rect 4433 15453 4445 15456
rect 4479 15453 4491 15487
rect 4433 15447 4491 15453
rect 4708 15487 4766 15493
rect 4708 15453 4720 15487
rect 4754 15453 4766 15487
rect 4708 15447 4766 15453
rect 4801 15487 4859 15493
rect 4801 15453 4813 15487
rect 4847 15484 4859 15487
rect 6181 15487 6239 15493
rect 6181 15484 6193 15487
rect 4847 15456 6193 15484
rect 4847 15453 4859 15456
rect 4801 15447 4859 15453
rect 6181 15453 6193 15456
rect 6227 15453 6239 15487
rect 6288 15484 6316 15592
rect 7006 15580 7012 15592
rect 7064 15580 7070 15632
rect 11606 15620 11612 15632
rect 11256 15592 11612 15620
rect 7466 15512 7472 15564
rect 7524 15552 7530 15564
rect 7837 15555 7895 15561
rect 7837 15552 7849 15555
rect 7524 15524 7849 15552
rect 7524 15512 7530 15524
rect 7837 15521 7849 15524
rect 7883 15552 7895 15555
rect 8021 15555 8079 15561
rect 8021 15552 8033 15555
rect 7883 15524 8033 15552
rect 7883 15521 7895 15524
rect 7837 15515 7895 15521
rect 8021 15521 8033 15524
rect 8067 15521 8079 15555
rect 8021 15515 8079 15521
rect 8481 15555 8539 15561
rect 8481 15521 8493 15555
rect 8527 15552 8539 15555
rect 9214 15552 9220 15564
rect 8527 15524 9220 15552
rect 8527 15521 8539 15524
rect 8481 15515 8539 15521
rect 9214 15512 9220 15524
rect 9272 15512 9278 15564
rect 11256 15561 11284 15592
rect 11606 15580 11612 15592
rect 11664 15580 11670 15632
rect 11716 15592 12388 15620
rect 10781 15555 10839 15561
rect 10781 15552 10793 15555
rect 9324 15524 10793 15552
rect 6365 15487 6423 15493
rect 6365 15484 6377 15487
rect 6288 15456 6377 15484
rect 6181 15447 6239 15453
rect 6365 15453 6377 15456
rect 6411 15453 6423 15487
rect 6365 15447 6423 15453
rect 6457 15487 6515 15493
rect 6457 15453 6469 15487
rect 6503 15453 6515 15487
rect 6457 15447 6515 15453
rect 2314 15376 2320 15428
rect 2372 15376 2378 15428
rect 2869 15419 2927 15425
rect 2869 15385 2881 15419
rect 2915 15385 2927 15419
rect 2869 15379 2927 15385
rect 3329 15419 3387 15425
rect 3329 15385 3341 15419
rect 3375 15416 3387 15419
rect 3375 15388 4476 15416
rect 3375 15385 3387 15388
rect 3329 15379 3387 15385
rect 2884 15348 2912 15379
rect 3789 15351 3847 15357
rect 3789 15348 3801 15351
rect 2884 15320 3801 15348
rect 3789 15317 3801 15320
rect 3835 15317 3847 15351
rect 4448 15348 4476 15388
rect 4816 15348 4844 15447
rect 6472 15416 6500 15447
rect 7650 15444 7656 15496
rect 7708 15493 7714 15496
rect 7708 15487 7725 15493
rect 7713 15486 7725 15487
rect 8389 15487 8447 15493
rect 7713 15484 7788 15486
rect 7713 15456 8340 15484
rect 7713 15453 7725 15456
rect 7708 15447 7725 15453
rect 7708 15444 7714 15447
rect 6825 15419 6883 15425
rect 6825 15416 6837 15419
rect 6472 15388 6837 15416
rect 6825 15385 6837 15388
rect 6871 15385 6883 15419
rect 6825 15379 6883 15385
rect 4448 15320 4844 15348
rect 6840 15348 6868 15379
rect 7006 15376 7012 15428
rect 7064 15376 7070 15428
rect 8312 15416 8340 15456
rect 8389 15453 8401 15487
rect 8435 15484 8447 15487
rect 9122 15484 9128 15496
rect 8435 15456 9128 15484
rect 8435 15453 8447 15456
rect 8389 15447 8447 15453
rect 9122 15444 9128 15456
rect 9180 15484 9186 15496
rect 9324 15484 9352 15524
rect 10781 15521 10793 15524
rect 10827 15521 10839 15555
rect 10781 15515 10839 15521
rect 11241 15555 11299 15561
rect 11241 15521 11253 15555
rect 11287 15521 11299 15555
rect 11716 15552 11744 15592
rect 11241 15515 11299 15521
rect 11440 15524 11744 15552
rect 12360 15552 12388 15592
rect 12618 15580 12624 15632
rect 12676 15620 12682 15632
rect 12676 15592 14504 15620
rect 12676 15580 12682 15592
rect 14090 15552 14096 15564
rect 12360 15524 14096 15552
rect 9180 15456 9352 15484
rect 9180 15444 9186 15456
rect 9582 15444 9588 15496
rect 9640 15444 9646 15496
rect 9950 15444 9956 15496
rect 10008 15444 10014 15496
rect 10045 15487 10103 15493
rect 10045 15453 10057 15487
rect 10091 15453 10103 15487
rect 10045 15447 10103 15453
rect 9769 15419 9827 15425
rect 9769 15416 9781 15419
rect 8312 15388 9781 15416
rect 9769 15385 9781 15388
rect 9815 15385 9827 15419
rect 10060 15416 10088 15447
rect 10410 15444 10416 15496
rect 10468 15484 10474 15496
rect 11440 15493 11468 15524
rect 14090 15512 14096 15524
rect 14148 15512 14154 15564
rect 14476 15561 14504 15592
rect 14918 15580 14924 15632
rect 14976 15580 14982 15632
rect 15102 15580 15108 15632
rect 15160 15620 15166 15632
rect 15197 15623 15255 15629
rect 15197 15620 15209 15623
rect 15160 15592 15209 15620
rect 15160 15580 15166 15592
rect 15197 15589 15209 15592
rect 15243 15589 15255 15623
rect 15197 15583 15255 15589
rect 14461 15555 14519 15561
rect 14461 15521 14473 15555
rect 14507 15552 14519 15555
rect 14550 15552 14556 15564
rect 14507 15524 14556 15552
rect 14507 15521 14519 15524
rect 14461 15515 14519 15521
rect 14550 15512 14556 15524
rect 14608 15512 14614 15564
rect 14936 15552 14964 15580
rect 15749 15555 15807 15561
rect 14660 15524 15424 15552
rect 10505 15487 10563 15493
rect 10505 15484 10517 15487
rect 10468 15456 10517 15484
rect 10468 15444 10474 15456
rect 10505 15453 10517 15456
rect 10551 15453 10563 15487
rect 10505 15447 10563 15453
rect 10689 15487 10747 15493
rect 10689 15453 10701 15487
rect 10735 15453 10747 15487
rect 10689 15447 10747 15453
rect 11149 15487 11207 15493
rect 11149 15453 11161 15487
rect 11195 15484 11207 15487
rect 11425 15487 11483 15493
rect 11425 15484 11437 15487
rect 11195 15456 11437 15484
rect 11195 15453 11207 15456
rect 11149 15447 11207 15453
rect 11425 15453 11437 15456
rect 11471 15453 11483 15487
rect 11425 15447 11483 15453
rect 10704 15416 10732 15447
rect 11606 15444 11612 15496
rect 11664 15444 11670 15496
rect 12161 15487 12219 15493
rect 12161 15453 12173 15487
rect 12207 15453 12219 15487
rect 12161 15447 12219 15453
rect 11238 15416 11244 15428
rect 10060 15388 11244 15416
rect 9769 15379 9827 15385
rect 11238 15376 11244 15388
rect 11296 15376 11302 15428
rect 6914 15348 6920 15360
rect 6840 15320 6920 15348
rect 3789 15311 3847 15317
rect 6914 15308 6920 15320
rect 6972 15348 6978 15360
rect 7469 15351 7527 15357
rect 7469 15348 7481 15351
rect 6972 15320 7481 15348
rect 6972 15308 6978 15320
rect 7469 15317 7481 15320
rect 7515 15317 7527 15351
rect 7469 15311 7527 15317
rect 8294 15308 8300 15360
rect 8352 15348 8358 15360
rect 8941 15351 8999 15357
rect 8941 15348 8953 15351
rect 8352 15320 8953 15348
rect 8352 15308 8358 15320
rect 8941 15317 8953 15320
rect 8987 15317 8999 15351
rect 8941 15311 8999 15317
rect 9125 15351 9183 15357
rect 9125 15317 9137 15351
rect 9171 15348 9183 15351
rect 9214 15348 9220 15360
rect 9171 15320 9220 15348
rect 9171 15317 9183 15320
rect 9125 15311 9183 15317
rect 9214 15308 9220 15320
rect 9272 15308 9278 15360
rect 10410 15308 10416 15360
rect 10468 15308 10474 15360
rect 10502 15308 10508 15360
rect 10560 15308 10566 15360
rect 12176 15348 12204 15447
rect 12342 15444 12348 15496
rect 12400 15444 12406 15496
rect 12434 15444 12440 15496
rect 12492 15444 12498 15496
rect 12529 15487 12587 15493
rect 12529 15453 12541 15487
rect 12575 15484 12587 15487
rect 12618 15484 12624 15496
rect 12575 15456 12624 15484
rect 12575 15453 12587 15456
rect 12529 15447 12587 15453
rect 12618 15444 12624 15456
rect 12676 15444 12682 15496
rect 12710 15444 12716 15496
rect 12768 15444 12774 15496
rect 12897 15487 12955 15493
rect 12897 15453 12909 15487
rect 12943 15484 12955 15487
rect 12989 15487 13047 15493
rect 12989 15484 13001 15487
rect 12943 15456 13001 15484
rect 12943 15453 12955 15456
rect 12897 15447 12955 15453
rect 12989 15453 13001 15456
rect 13035 15453 13047 15487
rect 12989 15447 13047 15453
rect 13354 15444 13360 15496
rect 13412 15444 13418 15496
rect 14660 15493 14688 15524
rect 14185 15487 14243 15493
rect 14185 15453 14197 15487
rect 14231 15453 14243 15487
rect 14185 15447 14243 15453
rect 14369 15487 14427 15493
rect 14369 15453 14381 15487
rect 14415 15484 14427 15487
rect 14645 15487 14703 15493
rect 14645 15484 14657 15487
rect 14415 15456 14657 15484
rect 14415 15453 14427 15456
rect 14369 15447 14427 15453
rect 14645 15453 14657 15456
rect 14691 15453 14703 15487
rect 14645 15447 14703 15453
rect 13170 15376 13176 15428
rect 13228 15376 13234 15428
rect 13265 15419 13323 15425
rect 13265 15385 13277 15419
rect 13311 15416 13323 15419
rect 13814 15416 13820 15428
rect 13311 15388 13820 15416
rect 13311 15385 13323 15388
rect 13265 15379 13323 15385
rect 13814 15376 13820 15388
rect 13872 15376 13878 15428
rect 14200 15416 14228 15447
rect 14826 15444 14832 15496
rect 14884 15444 14890 15496
rect 14918 15444 14924 15496
rect 14976 15444 14982 15496
rect 15102 15444 15108 15496
rect 15160 15444 15166 15496
rect 15396 15493 15424 15524
rect 15749 15521 15761 15555
rect 15795 15521 15807 15555
rect 15749 15515 15807 15521
rect 15197 15487 15255 15493
rect 15197 15453 15209 15487
rect 15243 15453 15255 15487
rect 15197 15447 15255 15453
rect 15381 15487 15439 15493
rect 15381 15453 15393 15487
rect 15427 15484 15439 15487
rect 15764 15484 15792 15515
rect 17218 15512 17224 15564
rect 17276 15512 17282 15564
rect 15427 15456 15792 15484
rect 15427 15453 15439 15456
rect 15381 15447 15439 15453
rect 14844 15416 14872 15444
rect 15212 15416 15240 15447
rect 17494 15444 17500 15496
rect 17552 15444 17558 15496
rect 15654 15416 15660 15428
rect 14200 15388 14412 15416
rect 14844 15388 15056 15416
rect 12526 15348 12532 15360
rect 12176 15320 12532 15348
rect 12526 15308 12532 15320
rect 12584 15308 12590 15360
rect 12710 15308 12716 15360
rect 12768 15348 12774 15360
rect 14277 15351 14335 15357
rect 14277 15348 14289 15351
rect 12768 15320 14289 15348
rect 12768 15308 12774 15320
rect 14277 15317 14289 15320
rect 14323 15317 14335 15351
rect 14384 15348 14412 15388
rect 14918 15348 14924 15360
rect 14384 15320 14924 15348
rect 14277 15311 14335 15317
rect 14918 15308 14924 15320
rect 14976 15308 14982 15360
rect 15028 15348 15056 15388
rect 15212 15388 15660 15416
rect 15212 15348 15240 15388
rect 15654 15376 15660 15388
rect 15712 15376 15718 15428
rect 16942 15416 16948 15428
rect 16790 15388 16948 15416
rect 16942 15376 16948 15388
rect 17000 15376 17006 15428
rect 15028 15320 15240 15348
rect 1104 15258 17848 15280
rect 1104 15206 2658 15258
rect 2710 15206 2722 15258
rect 2774 15206 2786 15258
rect 2838 15206 2850 15258
rect 2902 15206 2914 15258
rect 2966 15206 2978 15258
rect 3030 15206 8658 15258
rect 8710 15206 8722 15258
rect 8774 15206 8786 15258
rect 8838 15206 8850 15258
rect 8902 15206 8914 15258
rect 8966 15206 8978 15258
rect 9030 15206 14658 15258
rect 14710 15206 14722 15258
rect 14774 15206 14786 15258
rect 14838 15206 14850 15258
rect 14902 15206 14914 15258
rect 14966 15206 14978 15258
rect 15030 15206 17848 15258
rect 1104 15184 17848 15206
rect 1397 15147 1455 15153
rect 1397 15113 1409 15147
rect 1443 15144 1455 15147
rect 1578 15144 1584 15156
rect 1443 15116 1584 15144
rect 1443 15113 1455 15116
rect 1397 15107 1455 15113
rect 1578 15104 1584 15116
rect 1636 15104 1642 15156
rect 4246 15104 4252 15156
rect 4304 15104 4310 15156
rect 7834 15104 7840 15156
rect 7892 15144 7898 15156
rect 8021 15147 8079 15153
rect 8021 15144 8033 15147
rect 7892 15116 8033 15144
rect 7892 15104 7898 15116
rect 8021 15113 8033 15116
rect 8067 15113 8079 15147
rect 8021 15107 8079 15113
rect 8481 15147 8539 15153
rect 8481 15113 8493 15147
rect 8527 15113 8539 15147
rect 8481 15107 8539 15113
rect 8649 15147 8707 15153
rect 8649 15113 8661 15147
rect 8695 15144 8707 15147
rect 9582 15144 9588 15156
rect 8695 15116 9588 15144
rect 8695 15113 8707 15116
rect 8649 15107 8707 15113
rect 2406 15036 2412 15088
rect 2464 15036 2470 15088
rect 6914 15036 6920 15088
rect 6972 15036 6978 15088
rect 7101 15079 7159 15085
rect 7101 15045 7113 15079
rect 7147 15076 7159 15079
rect 7561 15079 7619 15085
rect 7561 15076 7573 15079
rect 7147 15048 7573 15076
rect 7147 15045 7159 15048
rect 7101 15039 7159 15045
rect 7561 15045 7573 15048
rect 7607 15045 7619 15079
rect 7561 15039 7619 15045
rect 7742 15036 7748 15088
rect 7800 15076 7806 15088
rect 8496 15076 8524 15107
rect 9582 15104 9588 15116
rect 9640 15104 9646 15156
rect 10410 15104 10416 15156
rect 10468 15144 10474 15156
rect 10689 15147 10747 15153
rect 10689 15144 10701 15147
rect 10468 15116 10701 15144
rect 10468 15104 10474 15116
rect 10689 15113 10701 15116
rect 10735 15113 10747 15147
rect 10689 15107 10747 15113
rect 12526 15104 12532 15156
rect 12584 15104 12590 15156
rect 12897 15147 12955 15153
rect 12897 15113 12909 15147
rect 12943 15144 12955 15147
rect 13170 15144 13176 15156
rect 12943 15116 13176 15144
rect 12943 15113 12955 15116
rect 12897 15107 12955 15113
rect 13170 15104 13176 15116
rect 13228 15104 13234 15156
rect 13909 15147 13967 15153
rect 13909 15113 13921 15147
rect 13955 15144 13967 15147
rect 14366 15144 14372 15156
rect 13955 15116 14372 15144
rect 13955 15113 13967 15116
rect 13909 15107 13967 15113
rect 14366 15104 14372 15116
rect 14424 15104 14430 15156
rect 15286 15104 15292 15156
rect 15344 15144 15350 15156
rect 16025 15147 16083 15153
rect 16025 15144 16037 15147
rect 15344 15116 16037 15144
rect 15344 15104 15350 15116
rect 16025 15113 16037 15116
rect 16071 15113 16083 15147
rect 16025 15107 16083 15113
rect 7800 15048 8524 15076
rect 8849 15079 8907 15085
rect 7800 15036 7806 15048
rect 4062 14968 4068 15020
rect 4120 15008 4126 15020
rect 4525 15011 4583 15017
rect 4525 15008 4537 15011
rect 4120 14980 4537 15008
rect 4120 14968 4126 14980
rect 4525 14977 4537 14980
rect 4571 14977 4583 15011
rect 4525 14971 4583 14977
rect 7466 14968 7472 15020
rect 7524 14968 7530 15020
rect 7650 14968 7656 15020
rect 7708 14968 7714 15020
rect 7852 15017 7880 15048
rect 8849 15045 8861 15079
rect 8895 15076 8907 15079
rect 9122 15076 9128 15088
rect 8895 15048 9128 15076
rect 8895 15045 8907 15048
rect 8849 15039 8907 15045
rect 9122 15036 9128 15048
rect 9180 15036 9186 15088
rect 10502 15076 10508 15088
rect 10152 15048 10508 15076
rect 7837 15011 7895 15017
rect 7837 14977 7849 15011
rect 7883 14977 7895 15011
rect 7837 14971 7895 14977
rect 8113 15011 8171 15017
rect 8113 14977 8125 15011
rect 8159 15008 8171 15011
rect 8294 15008 8300 15020
rect 8159 14980 8300 15008
rect 8159 14977 8171 14980
rect 8113 14971 8171 14977
rect 8294 14968 8300 14980
rect 8352 14968 8358 15020
rect 10152 15017 10180 15048
rect 10502 15036 10508 15048
rect 10560 15036 10566 15088
rect 12544 15076 12572 15104
rect 13630 15076 13636 15088
rect 12452 15048 13636 15076
rect 10137 15011 10195 15017
rect 10137 14977 10149 15011
rect 10183 14977 10195 15011
rect 10137 14971 10195 14977
rect 10413 15011 10471 15017
rect 10413 14977 10425 15011
rect 10459 15008 10471 15011
rect 11146 15008 11152 15020
rect 10459 14980 11152 15008
rect 10459 14977 10471 14980
rect 10413 14971 10471 14977
rect 11146 14968 11152 14980
rect 11204 14968 11210 15020
rect 12158 14968 12164 15020
rect 12216 14968 12222 15020
rect 12452 15017 12480 15048
rect 13630 15036 13636 15048
rect 13688 15036 13694 15088
rect 14458 15036 14464 15088
rect 14516 15076 14522 15088
rect 15013 15079 15071 15085
rect 14516 15048 14780 15076
rect 14516 15036 14522 15048
rect 12437 15011 12495 15017
rect 12437 14977 12449 15011
rect 12483 14977 12495 15011
rect 12437 14971 12495 14977
rect 12621 15011 12679 15017
rect 12621 14977 12633 15011
rect 12667 14977 12679 15011
rect 12621 14971 12679 14977
rect 2866 14900 2872 14952
rect 2924 14900 2930 14952
rect 3142 14900 3148 14952
rect 3200 14900 3206 14952
rect 4430 14900 4436 14952
rect 4488 14900 4494 14952
rect 4614 14900 4620 14952
rect 4672 14900 4678 14952
rect 4709 14943 4767 14949
rect 4709 14909 4721 14943
rect 4755 14940 4767 14943
rect 5350 14940 5356 14952
rect 4755 14912 5356 14940
rect 4755 14909 4767 14912
rect 4709 14903 4767 14909
rect 5350 14900 5356 14912
rect 5408 14900 5414 14952
rect 9950 14900 9956 14952
rect 10008 14940 10014 14952
rect 10229 14943 10287 14949
rect 10229 14940 10241 14943
rect 10008 14912 10241 14940
rect 10008 14900 10014 14912
rect 10229 14909 10241 14912
rect 10275 14909 10287 14943
rect 10229 14903 10287 14909
rect 10689 14943 10747 14949
rect 10689 14909 10701 14943
rect 10735 14940 10747 14943
rect 10870 14940 10876 14952
rect 10735 14912 10876 14940
rect 10735 14909 10747 14912
rect 10689 14903 10747 14909
rect 7006 14832 7012 14884
rect 7064 14872 7070 14884
rect 7837 14875 7895 14881
rect 7837 14872 7849 14875
rect 7064 14844 7849 14872
rect 7064 14832 7070 14844
rect 7837 14841 7849 14844
rect 7883 14841 7895 14875
rect 10244 14872 10272 14903
rect 10870 14900 10876 14912
rect 10928 14900 10934 14952
rect 11977 14875 12035 14881
rect 11977 14872 11989 14875
rect 10244 14844 11989 14872
rect 7837 14835 7895 14841
rect 11977 14841 11989 14844
rect 12023 14841 12035 14875
rect 12636 14872 12664 14971
rect 12710 14968 12716 15020
rect 12768 14968 12774 15020
rect 12802 14968 12808 15020
rect 12860 15008 12866 15020
rect 12897 15011 12955 15017
rect 12897 15008 12909 15011
rect 12860 14980 12909 15008
rect 12860 14968 12866 14980
rect 12897 14977 12909 14980
rect 12943 14977 12955 15011
rect 12897 14971 12955 14977
rect 13817 15011 13875 15017
rect 13817 14977 13829 15011
rect 13863 14977 13875 15011
rect 13817 14971 13875 14977
rect 14093 15011 14151 15017
rect 14093 14977 14105 15011
rect 14139 15008 14151 15011
rect 14185 15011 14243 15017
rect 14185 15008 14197 15011
rect 14139 14980 14197 15008
rect 14139 14977 14151 14980
rect 14093 14971 14151 14977
rect 14185 14977 14197 14980
rect 14231 14977 14243 15011
rect 14185 14971 14243 14977
rect 14369 15011 14427 15017
rect 14369 14977 14381 15011
rect 14415 14977 14427 15011
rect 14369 14971 14427 14977
rect 13170 14900 13176 14952
rect 13228 14940 13234 14952
rect 13354 14940 13360 14952
rect 13228 14912 13360 14940
rect 13228 14900 13234 14912
rect 13354 14900 13360 14912
rect 13412 14940 13418 14952
rect 13832 14940 13860 14971
rect 14384 14940 14412 14971
rect 14550 14968 14556 15020
rect 14608 14968 14614 15020
rect 14752 15017 14780 15048
rect 15013 15045 15025 15079
rect 15059 15045 15071 15079
rect 15013 15039 15071 15045
rect 14737 15011 14795 15017
rect 14737 14977 14749 15011
rect 14783 14977 14795 15011
rect 14737 14971 14795 14977
rect 14921 15011 14979 15017
rect 14921 14977 14933 15011
rect 14967 15008 14979 15011
rect 15028 15008 15056 15039
rect 14967 14980 15056 15008
rect 15289 15011 15347 15017
rect 14967 14977 14979 14980
rect 14921 14971 14979 14977
rect 15289 14977 15301 15011
rect 15335 15008 15347 15011
rect 15378 15008 15384 15020
rect 15335 14980 15384 15008
rect 15335 14977 15347 14980
rect 15289 14971 15347 14977
rect 13412 14912 13860 14940
rect 13924 14912 14412 14940
rect 13412 14900 13418 14912
rect 13078 14872 13084 14884
rect 12636 14844 13084 14872
rect 11977 14835 12035 14841
rect 13078 14832 13084 14844
rect 13136 14872 13142 14884
rect 13924 14872 13952 14912
rect 13136 14844 13952 14872
rect 13136 14832 13142 14844
rect 14090 14832 14096 14884
rect 14148 14832 14154 14884
rect 14384 14872 14412 14912
rect 14642 14900 14648 14952
rect 14700 14900 14706 14952
rect 15013 14943 15071 14949
rect 15013 14909 15025 14943
rect 15059 14940 15071 14943
rect 15102 14940 15108 14952
rect 15059 14912 15108 14940
rect 15059 14909 15071 14912
rect 15013 14903 15071 14909
rect 15102 14900 15108 14912
rect 15160 14900 15166 14952
rect 15304 14872 15332 14971
rect 15378 14968 15384 14980
rect 15436 14968 15442 15020
rect 15654 14968 15660 15020
rect 15712 14968 15718 15020
rect 16669 15011 16727 15017
rect 16669 14977 16681 15011
rect 16715 15008 16727 15011
rect 16758 15008 16764 15020
rect 16715 14980 16764 15008
rect 16715 14977 16727 14980
rect 16669 14971 16727 14977
rect 16758 14968 16764 14980
rect 16816 14968 16822 15020
rect 14384 14844 15332 14872
rect 15930 14832 15936 14884
rect 15988 14872 15994 14884
rect 16209 14875 16267 14881
rect 16209 14872 16221 14875
rect 15988 14844 16221 14872
rect 15988 14832 15994 14844
rect 16209 14841 16221 14844
rect 16255 14841 16267 14875
rect 16209 14835 16267 14841
rect 6086 14764 6092 14816
rect 6144 14804 6150 14816
rect 6733 14807 6791 14813
rect 6733 14804 6745 14807
rect 6144 14776 6745 14804
rect 6144 14764 6150 14776
rect 6733 14773 6745 14776
rect 6779 14773 6791 14807
rect 6733 14767 6791 14773
rect 8662 14764 8668 14816
rect 8720 14764 8726 14816
rect 8754 14764 8760 14816
rect 8812 14804 8818 14816
rect 9769 14807 9827 14813
rect 9769 14804 9781 14807
rect 8812 14776 9781 14804
rect 8812 14764 8818 14776
rect 9769 14773 9781 14776
rect 9815 14773 9827 14807
rect 9769 14767 9827 14773
rect 10505 14807 10563 14813
rect 10505 14773 10517 14807
rect 10551 14804 10563 14807
rect 11054 14804 11060 14816
rect 10551 14776 11060 14804
rect 10551 14773 10563 14776
rect 10505 14767 10563 14773
rect 11054 14764 11060 14776
rect 11112 14764 11118 14816
rect 12802 14764 12808 14816
rect 12860 14804 12866 14816
rect 13722 14804 13728 14816
rect 12860 14776 13728 14804
rect 12860 14764 12866 14776
rect 13722 14764 13728 14776
rect 13780 14804 13786 14816
rect 14642 14804 14648 14816
rect 13780 14776 14648 14804
rect 13780 14764 13786 14776
rect 14642 14764 14648 14776
rect 14700 14804 14706 14816
rect 15102 14804 15108 14816
rect 14700 14776 15108 14804
rect 14700 14764 14706 14776
rect 15102 14764 15108 14776
rect 15160 14764 15166 14816
rect 15197 14807 15255 14813
rect 15197 14773 15209 14807
rect 15243 14804 15255 14807
rect 15286 14804 15292 14816
rect 15243 14776 15292 14804
rect 15243 14773 15255 14776
rect 15197 14767 15255 14773
rect 15286 14764 15292 14776
rect 15344 14764 15350 14816
rect 16022 14764 16028 14816
rect 16080 14764 16086 14816
rect 16666 14764 16672 14816
rect 16724 14804 16730 14816
rect 16761 14807 16819 14813
rect 16761 14804 16773 14807
rect 16724 14776 16773 14804
rect 16724 14764 16730 14776
rect 16761 14773 16773 14776
rect 16807 14773 16819 14807
rect 16761 14767 16819 14773
rect 1104 14714 17848 14736
rect 1104 14662 1918 14714
rect 1970 14662 1982 14714
rect 2034 14662 2046 14714
rect 2098 14662 2110 14714
rect 2162 14662 2174 14714
rect 2226 14662 2238 14714
rect 2290 14662 7918 14714
rect 7970 14662 7982 14714
rect 8034 14662 8046 14714
rect 8098 14662 8110 14714
rect 8162 14662 8174 14714
rect 8226 14662 8238 14714
rect 8290 14662 13918 14714
rect 13970 14662 13982 14714
rect 14034 14662 14046 14714
rect 14098 14662 14110 14714
rect 14162 14662 14174 14714
rect 14226 14662 14238 14714
rect 14290 14662 17848 14714
rect 1104 14640 17848 14662
rect 2406 14560 2412 14612
rect 2464 14560 2470 14612
rect 2866 14560 2872 14612
rect 2924 14600 2930 14612
rect 3973 14603 4031 14609
rect 3973 14600 3985 14603
rect 2924 14572 3985 14600
rect 2924 14560 2930 14572
rect 3973 14569 3985 14572
rect 4019 14569 4031 14603
rect 3973 14563 4031 14569
rect 4338 14560 4344 14612
rect 4396 14600 4402 14612
rect 4433 14603 4491 14609
rect 4433 14600 4445 14603
rect 4396 14572 4445 14600
rect 4396 14560 4402 14572
rect 4433 14569 4445 14572
rect 4479 14569 4491 14603
rect 4433 14563 4491 14569
rect 5350 14560 5356 14612
rect 5408 14600 5414 14612
rect 5629 14603 5687 14609
rect 5629 14600 5641 14603
rect 5408 14572 5641 14600
rect 5408 14560 5414 14572
rect 5629 14569 5641 14572
rect 5675 14569 5687 14603
rect 5629 14563 5687 14569
rect 8662 14560 8668 14612
rect 8720 14600 8726 14612
rect 9214 14600 9220 14612
rect 8720 14572 9220 14600
rect 8720 14560 8726 14572
rect 9214 14560 9220 14572
rect 9272 14600 9278 14612
rect 9953 14603 10011 14609
rect 9953 14600 9965 14603
rect 9272 14572 9965 14600
rect 9272 14560 9278 14572
rect 9953 14569 9965 14572
rect 9999 14569 10011 14603
rect 9953 14563 10011 14569
rect 10870 14560 10876 14612
rect 10928 14560 10934 14612
rect 11054 14560 11060 14612
rect 11112 14560 11118 14612
rect 11238 14560 11244 14612
rect 11296 14600 11302 14612
rect 11425 14603 11483 14609
rect 11425 14600 11437 14603
rect 11296 14572 11437 14600
rect 11296 14560 11302 14572
rect 11425 14569 11437 14572
rect 11471 14569 11483 14603
rect 11425 14563 11483 14569
rect 12250 14560 12256 14612
rect 12308 14600 12314 14612
rect 13354 14600 13360 14612
rect 12308 14572 13360 14600
rect 12308 14560 12314 14572
rect 13354 14560 13360 14572
rect 13412 14560 13418 14612
rect 4709 14535 4767 14541
rect 4709 14501 4721 14535
rect 4755 14501 4767 14535
rect 6086 14532 6092 14544
rect 4709 14495 4767 14501
rect 5644 14504 6092 14532
rect 4724 14464 4752 14495
rect 3988 14436 4752 14464
rect 1394 14356 1400 14408
rect 1452 14396 1458 14408
rect 1581 14399 1639 14405
rect 1581 14396 1593 14399
rect 1452 14368 1593 14396
rect 1452 14356 1458 14368
rect 1581 14365 1593 14368
rect 1627 14365 1639 14399
rect 1581 14359 1639 14365
rect 2498 14356 2504 14408
rect 2556 14356 2562 14408
rect 3988 14405 4016 14436
rect 3973 14399 4031 14405
rect 3973 14365 3985 14399
rect 4019 14365 4031 14399
rect 3973 14359 4031 14365
rect 4154 14356 4160 14408
rect 4212 14356 4218 14408
rect 4982 14396 4988 14408
rect 4540 14368 4988 14396
rect 4062 14288 4068 14340
rect 4120 14328 4126 14340
rect 4430 14337 4436 14340
rect 4417 14331 4436 14337
rect 4120 14300 4384 14328
rect 4120 14288 4126 14300
rect 842 14220 848 14272
rect 900 14260 906 14272
rect 1397 14263 1455 14269
rect 1397 14260 1409 14263
rect 900 14232 1409 14260
rect 900 14220 906 14232
rect 1397 14229 1409 14232
rect 1443 14229 1455 14263
rect 1397 14223 1455 14229
rect 4154 14220 4160 14272
rect 4212 14260 4218 14272
rect 4249 14263 4307 14269
rect 4249 14260 4261 14263
rect 4212 14232 4261 14260
rect 4212 14220 4218 14232
rect 4249 14229 4261 14232
rect 4295 14229 4307 14263
rect 4356 14260 4384 14300
rect 4417 14297 4429 14331
rect 4488 14328 4494 14340
rect 4540 14328 4568 14368
rect 4982 14356 4988 14368
rect 5040 14356 5046 14408
rect 5350 14356 5356 14408
rect 5408 14356 5414 14408
rect 5644 14405 5672 14504
rect 6086 14492 6092 14504
rect 6144 14492 6150 14544
rect 5828 14436 6316 14464
rect 5828 14405 5856 14436
rect 5537 14399 5595 14405
rect 5537 14365 5549 14399
rect 5583 14365 5595 14399
rect 5537 14359 5595 14365
rect 5629 14399 5687 14405
rect 5629 14365 5641 14399
rect 5675 14365 5687 14399
rect 5629 14359 5687 14365
rect 5813 14399 5871 14405
rect 5813 14365 5825 14399
rect 5859 14365 5871 14399
rect 5813 14359 5871 14365
rect 4488 14300 4568 14328
rect 4417 14291 4436 14297
rect 4430 14288 4436 14291
rect 4488 14288 4494 14300
rect 4614 14288 4620 14340
rect 4672 14328 4678 14340
rect 4709 14331 4767 14337
rect 4709 14328 4721 14331
rect 4672 14300 4721 14328
rect 4672 14288 4678 14300
rect 4709 14297 4721 14300
rect 4755 14328 4767 14331
rect 5445 14331 5503 14337
rect 5445 14328 5457 14331
rect 4755 14300 5457 14328
rect 4755 14297 4767 14300
rect 4709 14291 4767 14297
rect 5445 14297 5457 14300
rect 5491 14297 5503 14331
rect 5552 14328 5580 14359
rect 6086 14356 6092 14408
rect 6144 14356 6150 14408
rect 6288 14405 6316 14436
rect 9858 14424 9864 14476
rect 9916 14464 9922 14476
rect 10505 14467 10563 14473
rect 10505 14464 10517 14467
rect 9916 14436 10517 14464
rect 9916 14424 9922 14436
rect 10505 14433 10517 14436
rect 10551 14464 10563 14467
rect 13814 14464 13820 14476
rect 10551 14436 13820 14464
rect 10551 14433 10563 14436
rect 10505 14427 10563 14433
rect 13814 14424 13820 14436
rect 13872 14424 13878 14476
rect 17494 14464 17500 14476
rect 15672 14436 17500 14464
rect 6273 14399 6331 14405
rect 6273 14365 6285 14399
rect 6319 14396 6331 14399
rect 6365 14399 6423 14405
rect 6365 14396 6377 14399
rect 6319 14368 6377 14396
rect 6319 14365 6331 14368
rect 6273 14359 6331 14365
rect 6365 14365 6377 14368
rect 6411 14365 6423 14399
rect 6365 14359 6423 14365
rect 6640 14399 6698 14405
rect 6640 14365 6652 14399
rect 6686 14365 6698 14399
rect 6640 14359 6698 14365
rect 6733 14399 6791 14405
rect 6733 14365 6745 14399
rect 6779 14396 6791 14399
rect 6822 14396 6828 14408
rect 6779 14368 6828 14396
rect 6779 14365 6791 14368
rect 6733 14359 6791 14365
rect 5905 14331 5963 14337
rect 5905 14328 5917 14331
rect 5552 14300 5917 14328
rect 5445 14291 5503 14297
rect 5905 14297 5917 14300
rect 5951 14297 5963 14331
rect 6656 14328 6684 14359
rect 6822 14356 6828 14368
rect 6880 14396 6886 14408
rect 8754 14396 8760 14408
rect 6880 14368 8760 14396
rect 6880 14356 6886 14368
rect 8754 14356 8760 14368
rect 8812 14356 8818 14408
rect 9766 14356 9772 14408
rect 9824 14396 9830 14408
rect 9953 14399 10011 14405
rect 9953 14396 9965 14399
rect 9824 14368 9965 14396
rect 9824 14356 9830 14368
rect 9953 14365 9965 14368
rect 9999 14365 10011 14399
rect 9953 14359 10011 14365
rect 10137 14399 10195 14405
rect 10137 14365 10149 14399
rect 10183 14365 10195 14399
rect 10137 14359 10195 14365
rect 10597 14399 10655 14405
rect 10597 14365 10609 14399
rect 10643 14396 10655 14399
rect 10686 14396 10692 14408
rect 10643 14368 10692 14396
rect 10643 14365 10655 14368
rect 10597 14359 10655 14365
rect 6914 14328 6920 14340
rect 6656 14300 6920 14328
rect 5905 14291 5963 14297
rect 6914 14288 6920 14300
rect 6972 14288 6978 14340
rect 10152 14328 10180 14359
rect 10686 14356 10692 14368
rect 10744 14356 10750 14408
rect 10870 14356 10876 14408
rect 10928 14396 10934 14408
rect 11057 14399 11115 14405
rect 11057 14396 11069 14399
rect 10928 14368 11069 14396
rect 10928 14356 10934 14368
rect 11057 14365 11069 14368
rect 11103 14365 11115 14399
rect 11057 14359 11115 14365
rect 11146 14356 11152 14408
rect 11204 14356 11210 14408
rect 13538 14356 13544 14408
rect 13596 14396 13602 14408
rect 15672 14405 15700 14436
rect 17494 14424 17500 14436
rect 17552 14424 17558 14476
rect 15657 14399 15715 14405
rect 15657 14396 15669 14399
rect 13596 14368 15669 14396
rect 13596 14356 13602 14368
rect 15657 14365 15669 14368
rect 15703 14365 15715 14399
rect 15657 14359 15715 14365
rect 11164 14328 11192 14356
rect 10152 14300 11192 14328
rect 15470 14288 15476 14340
rect 15528 14328 15534 14340
rect 15933 14331 15991 14337
rect 15933 14328 15945 14331
rect 15528 14300 15945 14328
rect 15528 14288 15534 14300
rect 15933 14297 15945 14300
rect 15979 14297 15991 14331
rect 15933 14291 15991 14297
rect 16666 14288 16672 14340
rect 16724 14288 16730 14340
rect 4893 14263 4951 14269
rect 4893 14260 4905 14263
rect 4356 14232 4905 14260
rect 4249 14223 4307 14229
rect 4893 14229 4905 14232
rect 4939 14229 4951 14263
rect 4893 14223 4951 14229
rect 17402 14220 17408 14272
rect 17460 14220 17466 14272
rect 1104 14170 17848 14192
rect 1104 14118 2658 14170
rect 2710 14118 2722 14170
rect 2774 14118 2786 14170
rect 2838 14118 2850 14170
rect 2902 14118 2914 14170
rect 2966 14118 2978 14170
rect 3030 14118 8658 14170
rect 8710 14118 8722 14170
rect 8774 14118 8786 14170
rect 8838 14118 8850 14170
rect 8902 14118 8914 14170
rect 8966 14118 8978 14170
rect 9030 14118 14658 14170
rect 14710 14118 14722 14170
rect 14774 14118 14786 14170
rect 14838 14118 14850 14170
rect 14902 14118 14914 14170
rect 14966 14118 14978 14170
rect 15030 14118 17848 14170
rect 1104 14096 17848 14118
rect 1394 14016 1400 14068
rect 1452 14016 1458 14068
rect 9766 14016 9772 14068
rect 9824 14016 9830 14068
rect 10962 14056 10968 14068
rect 9968 14028 10968 14056
rect 2314 13948 2320 14000
rect 2372 13948 2378 14000
rect 6733 13923 6791 13929
rect 6733 13889 6745 13923
rect 6779 13920 6791 13923
rect 6914 13920 6920 13932
rect 6779 13892 6920 13920
rect 6779 13889 6791 13892
rect 6733 13883 6791 13889
rect 6914 13880 6920 13892
rect 6972 13880 6978 13932
rect 9125 13923 9183 13929
rect 9125 13889 9137 13923
rect 9171 13920 9183 13923
rect 9490 13920 9496 13932
rect 9171 13892 9496 13920
rect 9171 13889 9183 13892
rect 9125 13883 9183 13889
rect 9490 13880 9496 13892
rect 9548 13880 9554 13932
rect 9677 13923 9735 13929
rect 9677 13889 9689 13923
rect 9723 13889 9735 13923
rect 9677 13883 9735 13889
rect 2866 13812 2872 13864
rect 2924 13812 2930 13864
rect 3142 13812 3148 13864
rect 3200 13812 3206 13864
rect 6822 13812 6828 13864
rect 6880 13812 6886 13864
rect 9306 13812 9312 13864
rect 9364 13812 9370 13864
rect 9407 13855 9465 13861
rect 9407 13821 9419 13855
rect 9453 13852 9465 13855
rect 9692 13852 9720 13883
rect 9858 13880 9864 13932
rect 9916 13880 9922 13932
rect 9968 13929 9996 14028
rect 10962 14016 10968 14028
rect 11020 14016 11026 14068
rect 11054 14016 11060 14068
rect 11112 14056 11118 14068
rect 11149 14059 11207 14065
rect 11149 14056 11161 14059
rect 11112 14028 11161 14056
rect 11112 14016 11118 14028
rect 11149 14025 11161 14028
rect 11195 14025 11207 14059
rect 11149 14019 11207 14025
rect 11606 14016 11612 14068
rect 11664 14056 11670 14068
rect 12253 14059 12311 14065
rect 12253 14056 12265 14059
rect 11664 14028 12265 14056
rect 11664 14016 11670 14028
rect 12253 14025 12265 14028
rect 12299 14025 12311 14059
rect 12253 14019 12311 14025
rect 12621 14059 12679 14065
rect 12621 14025 12633 14059
rect 12667 14056 12679 14059
rect 13262 14056 13268 14068
rect 12667 14028 13268 14056
rect 12667 14025 12679 14028
rect 12621 14019 12679 14025
rect 13262 14016 13268 14028
rect 13320 14016 13326 14068
rect 13446 14016 13452 14068
rect 13504 14016 13510 14068
rect 14277 14059 14335 14065
rect 14277 14025 14289 14059
rect 14323 14056 14335 14059
rect 14366 14056 14372 14068
rect 14323 14028 14372 14056
rect 14323 14025 14335 14028
rect 14277 14019 14335 14025
rect 14366 14016 14372 14028
rect 14424 14056 14430 14068
rect 14553 14059 14611 14065
rect 14553 14056 14565 14059
rect 14424 14028 14565 14056
rect 14424 14016 14430 14028
rect 14553 14025 14565 14028
rect 14599 14025 14611 14059
rect 15746 14056 15752 14068
rect 14553 14019 14611 14025
rect 14936 14028 15752 14056
rect 10045 13991 10103 13997
rect 10045 13957 10057 13991
rect 10091 13988 10103 13991
rect 12713 13991 12771 13997
rect 10091 13960 11100 13988
rect 10091 13957 10103 13960
rect 10045 13951 10103 13957
rect 9953 13923 10011 13929
rect 9953 13889 9965 13923
rect 9999 13889 10011 13923
rect 9953 13883 10011 13889
rect 10060 13852 10088 13951
rect 11072 13929 11100 13960
rect 12713 13957 12725 13991
rect 12759 13988 12771 13991
rect 14642 13988 14648 14000
rect 12759 13960 14648 13988
rect 12759 13957 12771 13960
rect 12713 13951 12771 13957
rect 14642 13948 14648 13960
rect 14700 13988 14706 14000
rect 14700 13960 14780 13988
rect 14700 13948 14706 13960
rect 10137 13923 10195 13929
rect 10137 13889 10149 13923
rect 10183 13889 10195 13923
rect 10137 13883 10195 13889
rect 10597 13923 10655 13929
rect 10597 13889 10609 13923
rect 10643 13920 10655 13923
rect 11057 13923 11115 13929
rect 10643 13892 11008 13920
rect 10643 13889 10655 13892
rect 10597 13883 10655 13889
rect 9453 13824 9536 13852
rect 9692 13824 10088 13852
rect 10152 13852 10180 13883
rect 10152 13824 10640 13852
rect 9453 13821 9465 13824
rect 9407 13815 9465 13821
rect 9508 13784 9536 13824
rect 9582 13784 9588 13796
rect 9508 13756 9588 13784
rect 9582 13744 9588 13756
rect 9640 13784 9646 13796
rect 10229 13787 10287 13793
rect 10229 13784 10241 13787
rect 9640 13756 10241 13784
rect 9640 13744 9646 13756
rect 10229 13753 10241 13756
rect 10275 13753 10287 13787
rect 10612 13784 10640 13824
rect 10686 13812 10692 13864
rect 10744 13812 10750 13864
rect 10980 13852 11008 13892
rect 11057 13889 11069 13923
rect 11103 13889 11115 13923
rect 11057 13883 11115 13889
rect 11238 13880 11244 13932
rect 11296 13880 11302 13932
rect 13078 13920 13084 13932
rect 12912 13892 13084 13920
rect 11256 13852 11284 13880
rect 12912 13861 12940 13892
rect 13078 13880 13084 13892
rect 13136 13880 13142 13932
rect 13354 13880 13360 13932
rect 13412 13880 13418 13932
rect 13722 13880 13728 13932
rect 13780 13920 13786 13932
rect 14752 13929 14780 13960
rect 14185 13923 14243 13929
rect 14185 13920 14197 13923
rect 13780 13892 14197 13920
rect 13780 13880 13786 13892
rect 14185 13889 14197 13892
rect 14231 13889 14243 13923
rect 14185 13883 14243 13889
rect 14461 13923 14519 13929
rect 14461 13889 14473 13923
rect 14507 13920 14519 13923
rect 14737 13923 14795 13929
rect 14507 13892 14688 13920
rect 14507 13889 14519 13892
rect 14461 13883 14519 13889
rect 10980 13824 11284 13852
rect 12897 13855 12955 13861
rect 12897 13821 12909 13855
rect 12943 13821 12955 13855
rect 12897 13815 12955 13821
rect 13173 13855 13231 13861
rect 13173 13821 13185 13855
rect 13219 13852 13231 13855
rect 13906 13852 13912 13864
rect 13219 13824 13912 13852
rect 13219 13821 13231 13824
rect 13173 13815 13231 13821
rect 11330 13784 11336 13796
rect 10612 13756 11336 13784
rect 10229 13747 10287 13753
rect 11330 13744 11336 13756
rect 11388 13744 11394 13796
rect 12342 13744 12348 13796
rect 12400 13784 12406 13796
rect 12526 13784 12532 13796
rect 12400 13756 12532 13784
rect 12400 13744 12406 13756
rect 12526 13744 12532 13756
rect 12584 13784 12590 13796
rect 12912 13784 12940 13815
rect 13906 13812 13912 13824
rect 13964 13852 13970 13864
rect 14660 13852 14688 13892
rect 14737 13889 14749 13923
rect 14783 13889 14795 13923
rect 14737 13883 14795 13889
rect 14936 13852 14964 14028
rect 15746 14016 15752 14028
rect 15804 14016 15810 14068
rect 16853 14059 16911 14065
rect 16853 14056 16865 14059
rect 15856 14028 16865 14056
rect 15013 13991 15071 13997
rect 15013 13957 15025 13991
rect 15059 13988 15071 13991
rect 15286 13988 15292 14000
rect 15059 13960 15292 13988
rect 15059 13957 15071 13960
rect 15013 13951 15071 13957
rect 15286 13948 15292 13960
rect 15344 13988 15350 14000
rect 15856 13997 15884 14028
rect 16853 14025 16865 14028
rect 16899 14025 16911 14059
rect 16853 14019 16911 14025
rect 15841 13991 15899 13997
rect 15841 13988 15853 13991
rect 15344 13960 15853 13988
rect 15344 13948 15350 13960
rect 15841 13957 15853 13960
rect 15887 13957 15899 13991
rect 15841 13951 15899 13957
rect 15102 13880 15108 13932
rect 15160 13920 15166 13932
rect 15197 13923 15255 13929
rect 15197 13920 15209 13923
rect 15160 13892 15209 13920
rect 15160 13880 15166 13892
rect 15197 13889 15209 13892
rect 15243 13920 15255 13923
rect 15243 13892 15332 13920
rect 15243 13889 15255 13892
rect 15197 13883 15255 13889
rect 13964 13824 14504 13852
rect 14660 13824 14964 13852
rect 13964 13812 13970 13824
rect 14476 13796 14504 13824
rect 12584 13756 12940 13784
rect 12584 13744 12590 13756
rect 14458 13744 14464 13796
rect 14516 13744 14522 13796
rect 15304 13784 15332 13892
rect 15378 13880 15384 13932
rect 15436 13920 15442 13932
rect 15657 13923 15715 13929
rect 15657 13920 15669 13923
rect 15436 13892 15669 13920
rect 15436 13880 15442 13892
rect 15657 13889 15669 13892
rect 15703 13920 15715 13923
rect 16022 13920 16028 13932
rect 15703 13892 16028 13920
rect 15703 13889 15715 13892
rect 15657 13883 15715 13889
rect 16022 13880 16028 13892
rect 16080 13880 16086 13932
rect 16850 13880 16856 13932
rect 16908 13920 16914 13932
rect 17037 13923 17095 13929
rect 17037 13920 17049 13923
rect 16908 13892 17049 13920
rect 16908 13880 16914 13892
rect 17037 13889 17049 13892
rect 17083 13889 17095 13923
rect 17037 13883 17095 13889
rect 16574 13812 16580 13864
rect 16632 13852 16638 13864
rect 16669 13855 16727 13861
rect 16669 13852 16681 13855
rect 16632 13824 16681 13852
rect 16632 13812 16638 13824
rect 16669 13821 16681 13824
rect 16715 13821 16727 13855
rect 16669 13815 16727 13821
rect 15654 13784 15660 13796
rect 15304 13756 15660 13784
rect 15654 13744 15660 13756
rect 15712 13744 15718 13796
rect 6362 13676 6368 13728
rect 6420 13716 6426 13728
rect 6457 13719 6515 13725
rect 6457 13716 6469 13719
rect 6420 13688 6469 13716
rect 6420 13676 6426 13688
rect 6457 13685 6469 13688
rect 6503 13685 6515 13719
rect 6457 13679 6515 13685
rect 8478 13676 8484 13728
rect 8536 13716 8542 13728
rect 8941 13719 8999 13725
rect 8941 13716 8953 13719
rect 8536 13688 8953 13716
rect 8536 13676 8542 13688
rect 8941 13685 8953 13688
rect 8987 13685 8999 13719
rect 8941 13679 8999 13685
rect 14918 13676 14924 13728
rect 14976 13676 14982 13728
rect 15378 13676 15384 13728
rect 15436 13676 15442 13728
rect 15470 13676 15476 13728
rect 15528 13676 15534 13728
rect 17221 13719 17279 13725
rect 17221 13685 17233 13719
rect 17267 13716 17279 13719
rect 17402 13716 17408 13728
rect 17267 13688 17408 13716
rect 17267 13685 17279 13688
rect 17221 13679 17279 13685
rect 17402 13676 17408 13688
rect 17460 13676 17466 13728
rect 1104 13626 17848 13648
rect 1104 13574 1918 13626
rect 1970 13574 1982 13626
rect 2034 13574 2046 13626
rect 2098 13574 2110 13626
rect 2162 13574 2174 13626
rect 2226 13574 2238 13626
rect 2290 13574 7918 13626
rect 7970 13574 7982 13626
rect 8034 13574 8046 13626
rect 8098 13574 8110 13626
rect 8162 13574 8174 13626
rect 8226 13574 8238 13626
rect 8290 13574 13918 13626
rect 13970 13574 13982 13626
rect 14034 13574 14046 13626
rect 14098 13574 14110 13626
rect 14162 13574 14174 13626
rect 14226 13574 14238 13626
rect 14290 13574 17848 13626
rect 1104 13552 17848 13574
rect 2314 13472 2320 13524
rect 2372 13472 2378 13524
rect 2866 13472 2872 13524
rect 2924 13512 2930 13524
rect 2961 13515 3019 13521
rect 2961 13512 2973 13515
rect 2924 13484 2973 13512
rect 2924 13472 2930 13484
rect 2961 13481 2973 13484
rect 3007 13481 3019 13515
rect 2961 13475 3019 13481
rect 5258 13472 5264 13524
rect 5316 13512 5322 13524
rect 5537 13515 5595 13521
rect 5537 13512 5549 13515
rect 5316 13484 5549 13512
rect 5316 13472 5322 13484
rect 5537 13481 5549 13484
rect 5583 13512 5595 13515
rect 6365 13515 6423 13521
rect 6365 13512 6377 13515
rect 5583 13484 6377 13512
rect 5583 13481 5595 13484
rect 5537 13475 5595 13481
rect 6365 13481 6377 13484
rect 6411 13481 6423 13515
rect 6365 13475 6423 13481
rect 7650 13472 7656 13524
rect 7708 13512 7714 13524
rect 8021 13515 8079 13521
rect 8021 13512 8033 13515
rect 7708 13484 8033 13512
rect 7708 13472 7714 13484
rect 8021 13481 8033 13484
rect 8067 13481 8079 13515
rect 8021 13475 8079 13481
rect 11146 13472 11152 13524
rect 11204 13472 11210 13524
rect 13262 13472 13268 13524
rect 13320 13512 13326 13524
rect 13906 13512 13912 13524
rect 13320 13484 13912 13512
rect 13320 13472 13326 13484
rect 13906 13472 13912 13484
rect 13964 13472 13970 13524
rect 6181 13447 6239 13453
rect 6181 13444 6193 13447
rect 5368 13416 6193 13444
rect 5368 13388 5396 13416
rect 6181 13413 6193 13416
rect 6227 13413 6239 13447
rect 6181 13407 6239 13413
rect 7929 13447 7987 13453
rect 7929 13413 7941 13447
rect 7975 13413 7987 13447
rect 7929 13407 7987 13413
rect 3329 13379 3387 13385
rect 3329 13345 3341 13379
rect 3375 13376 3387 13379
rect 4893 13379 4951 13385
rect 4893 13376 4905 13379
rect 3375 13348 4905 13376
rect 3375 13345 3387 13348
rect 3329 13339 3387 13345
rect 4893 13345 4905 13348
rect 4939 13345 4951 13379
rect 5350 13376 5356 13388
rect 4893 13339 4951 13345
rect 5184 13348 5356 13376
rect 1394 13268 1400 13320
rect 1452 13308 1458 13320
rect 1581 13311 1639 13317
rect 1581 13308 1593 13311
rect 1452 13280 1593 13308
rect 1452 13268 1458 13280
rect 1581 13277 1593 13280
rect 1627 13277 1639 13311
rect 1581 13271 1639 13277
rect 2409 13311 2467 13317
rect 2409 13277 2421 13311
rect 2455 13308 2467 13311
rect 2498 13308 2504 13320
rect 2455 13280 2504 13308
rect 2455 13277 2467 13280
rect 2409 13271 2467 13277
rect 2498 13268 2504 13280
rect 2556 13268 2562 13320
rect 3237 13311 3295 13317
rect 3237 13277 3249 13311
rect 3283 13308 3295 13311
rect 3510 13308 3516 13320
rect 3283 13280 3516 13308
rect 3283 13277 3295 13280
rect 3237 13271 3295 13277
rect 3510 13268 3516 13280
rect 3568 13268 3574 13320
rect 5184 13317 5212 13348
rect 5350 13336 5356 13348
rect 5408 13336 5414 13388
rect 7653 13379 7711 13385
rect 6104 13348 6592 13376
rect 5258 13317 5264 13320
rect 5168 13311 5226 13317
rect 5168 13277 5180 13311
rect 5214 13277 5226 13311
rect 5168 13271 5226 13277
rect 5254 13271 5264 13317
rect 5316 13308 5322 13320
rect 5316 13280 5354 13308
rect 5258 13268 5264 13271
rect 5316 13268 5322 13280
rect 5626 13268 5632 13320
rect 5684 13268 5690 13320
rect 6104 13317 6132 13348
rect 6089 13311 6147 13317
rect 6089 13277 6101 13311
rect 6135 13277 6147 13311
rect 6089 13271 6147 13277
rect 6273 13311 6331 13317
rect 6273 13277 6285 13311
rect 6319 13308 6331 13311
rect 6362 13308 6368 13320
rect 6319 13280 6368 13308
rect 6319 13277 6331 13280
rect 6273 13271 6331 13277
rect 6362 13268 6368 13280
rect 6420 13268 6426 13320
rect 6564 13317 6592 13348
rect 7653 13345 7665 13379
rect 7699 13376 7711 13379
rect 7742 13376 7748 13388
rect 7699 13348 7748 13376
rect 7699 13345 7711 13348
rect 7653 13339 7711 13345
rect 7742 13336 7748 13348
rect 7800 13336 7806 13388
rect 6549 13311 6607 13317
rect 6549 13277 6561 13311
rect 6595 13308 6607 13311
rect 7098 13308 7104 13320
rect 6595 13280 7104 13308
rect 6595 13277 6607 13280
rect 6549 13271 6607 13277
rect 7098 13268 7104 13280
rect 7156 13268 7162 13320
rect 7558 13268 7564 13320
rect 7616 13268 7622 13320
rect 7944 13308 7972 13407
rect 13814 13404 13820 13456
rect 13872 13444 13878 13456
rect 14185 13447 14243 13453
rect 14185 13444 14197 13447
rect 13872 13416 14197 13444
rect 13872 13404 13878 13416
rect 14185 13413 14197 13416
rect 14231 13413 14243 13447
rect 14185 13407 14243 13413
rect 14642 13404 14648 13456
rect 14700 13444 14706 13456
rect 14700 13416 16436 13444
rect 14700 13404 14706 13416
rect 16408 13388 16436 13416
rect 8481 13379 8539 13385
rect 8481 13345 8493 13379
rect 8527 13376 8539 13379
rect 9490 13376 9496 13388
rect 8527 13348 9496 13376
rect 8527 13345 8539 13348
rect 8481 13339 8539 13345
rect 9490 13336 9496 13348
rect 9548 13336 9554 13388
rect 11054 13336 11060 13388
rect 11112 13376 11118 13388
rect 11517 13379 11575 13385
rect 11517 13376 11529 13379
rect 11112 13348 11529 13376
rect 11112 13336 11118 13348
rect 11517 13345 11529 13348
rect 11563 13345 11575 13379
rect 11517 13339 11575 13345
rect 11974 13336 11980 13388
rect 12032 13376 12038 13388
rect 12802 13376 12808 13388
rect 12032 13348 12808 13376
rect 12032 13336 12038 13348
rect 12802 13336 12808 13348
rect 12860 13336 12866 13388
rect 14918 13336 14924 13388
rect 14976 13376 14982 13388
rect 14976 13348 15792 13376
rect 14976 13336 14982 13348
rect 8389 13311 8447 13317
rect 8389 13308 8401 13311
rect 7944 13280 8401 13308
rect 8389 13277 8401 13280
rect 8435 13277 8447 13311
rect 8389 13271 8447 13277
rect 8941 13311 8999 13317
rect 8941 13277 8953 13311
rect 8987 13308 8999 13311
rect 10134 13308 10140 13320
rect 8987 13280 10140 13308
rect 8987 13277 8999 13280
rect 8941 13271 8999 13277
rect 8956 13240 8984 13271
rect 10134 13268 10140 13280
rect 10192 13268 10198 13320
rect 11330 13268 11336 13320
rect 11388 13268 11394 13320
rect 11885 13311 11943 13317
rect 11885 13277 11897 13311
rect 11931 13308 11943 13311
rect 12158 13308 12164 13320
rect 11931 13280 12164 13308
rect 11931 13277 11943 13280
rect 11885 13271 11943 13277
rect 12158 13268 12164 13280
rect 12216 13308 12222 13320
rect 13538 13308 13544 13320
rect 12216 13280 13544 13308
rect 12216 13268 12222 13280
rect 13538 13268 13544 13280
rect 13596 13268 13602 13320
rect 14369 13311 14427 13317
rect 14369 13277 14381 13311
rect 14415 13308 14427 13311
rect 14458 13308 14464 13320
rect 14415 13280 14464 13308
rect 14415 13277 14427 13280
rect 14369 13271 14427 13277
rect 14458 13268 14464 13280
rect 14516 13268 14522 13320
rect 14734 13268 14740 13320
rect 14792 13268 14798 13320
rect 14829 13311 14887 13317
rect 14829 13277 14841 13311
rect 14875 13277 14887 13311
rect 14829 13271 14887 13277
rect 6380 13212 8984 13240
rect 6380 13184 6408 13212
rect 9674 13200 9680 13252
rect 9732 13240 9738 13252
rect 11977 13243 12035 13249
rect 11977 13240 11989 13243
rect 9732 13212 11989 13240
rect 9732 13200 9738 13212
rect 11977 13209 11989 13212
rect 12023 13209 12035 13243
rect 11977 13203 12035 13209
rect 14274 13200 14280 13252
rect 14332 13240 14338 13252
rect 14844 13240 14872 13271
rect 15378 13268 15384 13320
rect 15436 13268 15442 13320
rect 15764 13317 15792 13348
rect 16390 13336 16396 13388
rect 16448 13336 16454 13388
rect 17402 13376 17408 13388
rect 16776 13348 17408 13376
rect 16776 13320 16804 13348
rect 17402 13336 17408 13348
rect 17460 13336 17466 13388
rect 15749 13311 15807 13317
rect 15749 13277 15761 13311
rect 15795 13277 15807 13311
rect 15749 13271 15807 13277
rect 16209 13311 16267 13317
rect 16209 13277 16221 13311
rect 16255 13308 16267 13311
rect 16574 13308 16580 13320
rect 16255 13280 16580 13308
rect 16255 13277 16267 13280
rect 16209 13271 16267 13277
rect 16574 13268 16580 13280
rect 16632 13268 16638 13320
rect 16758 13268 16764 13320
rect 16816 13268 16822 13320
rect 16850 13268 16856 13320
rect 16908 13268 16914 13320
rect 14332 13212 14872 13240
rect 14332 13200 14338 13212
rect 842 13132 848 13184
rect 900 13172 906 13184
rect 1397 13175 1455 13181
rect 1397 13172 1409 13175
rect 900 13144 1409 13172
rect 900 13132 906 13144
rect 1397 13141 1409 13144
rect 1443 13141 1455 13175
rect 1397 13135 1455 13141
rect 4982 13132 4988 13184
rect 5040 13172 5046 13184
rect 5353 13175 5411 13181
rect 5353 13172 5365 13175
rect 5040 13144 5365 13172
rect 5040 13132 5046 13144
rect 5353 13141 5365 13144
rect 5399 13141 5411 13175
rect 5353 13135 5411 13141
rect 6362 13132 6368 13184
rect 6420 13132 6426 13184
rect 12066 13132 12072 13184
rect 12124 13172 12130 13184
rect 12710 13172 12716 13184
rect 12124 13144 12716 13172
rect 12124 13132 12130 13144
rect 12710 13132 12716 13144
rect 12768 13132 12774 13184
rect 13538 13132 13544 13184
rect 13596 13172 13602 13184
rect 13722 13172 13728 13184
rect 13596 13144 13728 13172
rect 13596 13132 13602 13144
rect 13722 13132 13728 13144
rect 13780 13132 13786 13184
rect 14458 13132 14464 13184
rect 14516 13172 14522 13184
rect 14734 13172 14740 13184
rect 14516 13144 14740 13172
rect 14516 13132 14522 13144
rect 14734 13132 14740 13144
rect 14792 13172 14798 13184
rect 16206 13172 16212 13184
rect 14792 13144 16212 13172
rect 14792 13132 14798 13144
rect 16206 13132 16212 13144
rect 16264 13132 16270 13184
rect 1104 13082 17848 13104
rect 1104 13030 2658 13082
rect 2710 13030 2722 13082
rect 2774 13030 2786 13082
rect 2838 13030 2850 13082
rect 2902 13030 2914 13082
rect 2966 13030 2978 13082
rect 3030 13030 8658 13082
rect 8710 13030 8722 13082
rect 8774 13030 8786 13082
rect 8838 13030 8850 13082
rect 8902 13030 8914 13082
rect 8966 13030 8978 13082
rect 9030 13030 14658 13082
rect 14710 13030 14722 13082
rect 14774 13030 14786 13082
rect 14838 13030 14850 13082
rect 14902 13030 14914 13082
rect 14966 13030 14978 13082
rect 15030 13030 17848 13082
rect 1104 13008 17848 13030
rect 1394 12928 1400 12980
rect 1452 12928 1458 12980
rect 3510 12928 3516 12980
rect 3568 12928 3574 12980
rect 5350 12928 5356 12980
rect 5408 12968 5414 12980
rect 5408 12940 5488 12968
rect 5408 12928 5414 12940
rect 2314 12860 2320 12912
rect 2372 12860 2378 12912
rect 3160 12872 5120 12900
rect 3160 12841 3188 12872
rect 3145 12835 3203 12841
rect 3145 12801 3157 12835
rect 3191 12801 3203 12835
rect 3145 12795 3203 12801
rect 3418 12792 3424 12844
rect 3476 12792 3482 12844
rect 3605 12835 3663 12841
rect 3605 12801 3617 12835
rect 3651 12832 3663 12835
rect 4706 12832 4712 12844
rect 4764 12841 4770 12844
rect 4764 12835 4797 12841
rect 3651 12804 4712 12832
rect 3651 12801 3663 12804
rect 3605 12795 3663 12801
rect 4706 12792 4712 12804
rect 4785 12801 4797 12835
rect 4764 12795 4797 12801
rect 4893 12835 4951 12841
rect 4893 12801 4905 12835
rect 4939 12801 4951 12835
rect 4893 12795 4951 12801
rect 4764 12792 4770 12795
rect 2869 12767 2927 12773
rect 2869 12733 2881 12767
rect 2915 12764 2927 12767
rect 2915 12736 3096 12764
rect 2915 12733 2927 12736
rect 2869 12727 2927 12733
rect 3068 12696 3096 12736
rect 3602 12696 3608 12708
rect 3068 12668 3608 12696
rect 3602 12656 3608 12668
rect 3660 12656 3666 12708
rect 4246 12656 4252 12708
rect 4304 12696 4310 12708
rect 4525 12699 4583 12705
rect 4525 12696 4537 12699
rect 4304 12668 4537 12696
rect 4304 12656 4310 12668
rect 4525 12665 4537 12668
rect 4571 12665 4583 12699
rect 4908 12696 4936 12795
rect 4982 12724 4988 12776
rect 5040 12724 5046 12776
rect 5092 12764 5120 12872
rect 5166 12792 5172 12844
rect 5224 12832 5230 12844
rect 5261 12835 5319 12841
rect 5261 12832 5273 12835
rect 5224 12804 5273 12832
rect 5224 12792 5230 12804
rect 5261 12801 5273 12804
rect 5307 12801 5319 12835
rect 5261 12795 5319 12801
rect 5350 12792 5356 12844
rect 5408 12792 5414 12844
rect 5460 12841 5488 12940
rect 7558 12928 7564 12980
rect 7616 12968 7622 12980
rect 8297 12971 8355 12977
rect 8297 12968 8309 12971
rect 7616 12940 8309 12968
rect 7616 12928 7622 12940
rect 8297 12937 8309 12940
rect 8343 12968 8355 12971
rect 9582 12968 9588 12980
rect 8343 12940 9588 12968
rect 8343 12937 8355 12940
rect 8297 12931 8355 12937
rect 9582 12928 9588 12940
rect 9640 12928 9646 12980
rect 10134 12928 10140 12980
rect 10192 12968 10198 12980
rect 11054 12968 11060 12980
rect 10192 12940 11060 12968
rect 10192 12928 10198 12940
rect 11054 12928 11060 12940
rect 11112 12928 11118 12980
rect 12434 12928 12440 12980
rect 12492 12968 12498 12980
rect 12894 12968 12900 12980
rect 12492 12940 12900 12968
rect 12492 12928 12498 12940
rect 12894 12928 12900 12940
rect 12952 12928 12958 12980
rect 13446 12928 13452 12980
rect 13504 12928 13510 12980
rect 14274 12928 14280 12980
rect 14332 12928 14338 12980
rect 14458 12928 14464 12980
rect 14516 12928 14522 12980
rect 15197 12971 15255 12977
rect 15197 12968 15209 12971
rect 14752 12940 15209 12968
rect 8113 12903 8171 12909
rect 8113 12869 8125 12903
rect 8159 12900 8171 12903
rect 8849 12903 8907 12909
rect 8849 12900 8861 12903
rect 8159 12872 8861 12900
rect 8159 12869 8171 12872
rect 8113 12863 8171 12869
rect 8849 12869 8861 12872
rect 8895 12900 8907 12903
rect 9674 12900 9680 12912
rect 8895 12872 9680 12900
rect 8895 12869 8907 12872
rect 8849 12863 8907 12869
rect 9674 12860 9680 12872
rect 9732 12860 9738 12912
rect 11146 12900 11152 12912
rect 11072 12872 11152 12900
rect 5445 12835 5503 12841
rect 5445 12801 5457 12835
rect 5491 12801 5503 12835
rect 5445 12795 5503 12801
rect 5534 12792 5540 12844
rect 5592 12832 5598 12844
rect 5629 12835 5687 12841
rect 5629 12832 5641 12835
rect 5592 12804 5641 12832
rect 5592 12792 5598 12804
rect 5629 12801 5641 12804
rect 5675 12801 5687 12835
rect 5629 12795 5687 12801
rect 7742 12792 7748 12844
rect 7800 12832 7806 12844
rect 8205 12835 8263 12841
rect 8205 12832 8217 12835
rect 7800 12804 8217 12832
rect 7800 12792 7806 12804
rect 8205 12801 8217 12804
rect 8251 12801 8263 12835
rect 8205 12795 8263 12801
rect 6362 12764 6368 12776
rect 5092 12736 6368 12764
rect 6362 12724 6368 12736
rect 6420 12724 6426 12776
rect 8220 12764 8248 12795
rect 8478 12792 8484 12844
rect 8536 12792 8542 12844
rect 11072 12841 11100 12872
rect 11146 12860 11152 12872
rect 11204 12900 11210 12912
rect 11606 12900 11612 12912
rect 11204 12872 11612 12900
rect 11204 12860 11210 12872
rect 11606 12860 11612 12872
rect 11664 12860 11670 12912
rect 12069 12903 12127 12909
rect 12069 12869 12081 12903
rect 12115 12900 12127 12903
rect 12115 12872 12296 12900
rect 12115 12869 12127 12872
rect 12069 12863 12127 12869
rect 11057 12835 11115 12841
rect 11057 12801 11069 12835
rect 11103 12801 11115 12835
rect 11057 12795 11115 12801
rect 11974 12792 11980 12844
rect 12032 12792 12038 12844
rect 12268 12841 12296 12872
rect 12452 12841 12480 12928
rect 13354 12900 13360 12912
rect 12544 12872 13360 12900
rect 12544 12841 12572 12872
rect 13354 12860 13360 12872
rect 13412 12860 13418 12912
rect 14476 12900 14504 12928
rect 14752 12909 14780 12940
rect 15197 12937 15209 12940
rect 15243 12937 15255 12971
rect 15197 12931 15255 12937
rect 16206 12928 16212 12980
rect 16264 12928 16270 12980
rect 14599 12903 14657 12909
rect 14599 12900 14611 12903
rect 14476 12872 14611 12900
rect 14599 12869 14611 12872
rect 14645 12869 14657 12903
rect 14599 12863 14657 12869
rect 14737 12903 14795 12909
rect 14737 12869 14749 12903
rect 14783 12869 14795 12903
rect 14737 12863 14795 12869
rect 14829 12903 14887 12909
rect 14829 12869 14841 12903
rect 14875 12900 14887 12903
rect 15470 12900 15476 12912
rect 14875 12872 15476 12900
rect 14875 12869 14887 12872
rect 14829 12863 14887 12869
rect 15470 12860 15476 12872
rect 15528 12860 15534 12912
rect 12161 12835 12219 12841
rect 12161 12801 12173 12835
rect 12207 12801 12219 12835
rect 12161 12795 12219 12801
rect 12253 12835 12311 12841
rect 12253 12801 12265 12835
rect 12299 12801 12311 12835
rect 12253 12795 12311 12801
rect 12437 12835 12495 12841
rect 12437 12801 12449 12835
rect 12483 12801 12495 12835
rect 12437 12795 12495 12801
rect 12529 12835 12587 12841
rect 12529 12801 12541 12835
rect 12575 12801 12587 12835
rect 12529 12795 12587 12801
rect 9306 12764 9312 12776
rect 8220 12736 9312 12764
rect 9306 12724 9312 12736
rect 9364 12724 9370 12776
rect 9490 12724 9496 12776
rect 9548 12764 9554 12776
rect 9548 12736 11100 12764
rect 9548 12724 9554 12736
rect 5626 12696 5632 12708
rect 4908 12668 5632 12696
rect 4525 12659 4583 12665
rect 5626 12656 5632 12668
rect 5684 12656 5690 12708
rect 6914 12656 6920 12708
rect 6972 12696 6978 12708
rect 8481 12699 8539 12705
rect 8481 12696 8493 12699
rect 6972 12668 8493 12696
rect 6972 12656 6978 12668
rect 8481 12665 8493 12668
rect 8527 12665 8539 12699
rect 8481 12659 8539 12665
rect 10686 12656 10692 12708
rect 10744 12656 10750 12708
rect 11072 12696 11100 12736
rect 11146 12724 11152 12776
rect 11204 12764 11210 12776
rect 11330 12764 11336 12776
rect 11204 12736 11336 12764
rect 11204 12724 11210 12736
rect 11330 12724 11336 12736
rect 11388 12724 11394 12776
rect 12066 12724 12072 12776
rect 12124 12764 12130 12776
rect 12176 12764 12204 12795
rect 12618 12792 12624 12844
rect 12676 12792 12682 12844
rect 12802 12792 12808 12844
rect 12860 12792 12866 12844
rect 13078 12792 13084 12844
rect 13136 12832 13142 12844
rect 13909 12835 13967 12841
rect 13136 12804 13768 12832
rect 13136 12792 13142 12804
rect 12989 12767 13047 12773
rect 12124 12736 12204 12764
rect 12268 12736 12664 12764
rect 12124 12724 12130 12736
rect 12268 12696 12296 12736
rect 11072 12668 12296 12696
rect 12636 12696 12664 12736
rect 12989 12733 13001 12767
rect 13035 12764 13047 12767
rect 13541 12767 13599 12773
rect 13541 12764 13553 12767
rect 13035 12736 13553 12764
rect 13035 12733 13047 12736
rect 12989 12727 13047 12733
rect 13541 12733 13553 12736
rect 13587 12733 13599 12767
rect 13541 12727 13599 12733
rect 13630 12724 13636 12776
rect 13688 12724 13694 12776
rect 13740 12764 13768 12804
rect 13909 12801 13921 12835
rect 13955 12832 13967 12835
rect 14274 12832 14280 12844
rect 13955 12804 14280 12832
rect 13955 12801 13967 12804
rect 13909 12795 13967 12801
rect 14274 12792 14280 12804
rect 14332 12792 14338 12844
rect 14366 12792 14372 12844
rect 14424 12832 14430 12844
rect 14461 12835 14519 12841
rect 14461 12832 14473 12835
rect 14424 12804 14473 12832
rect 14424 12792 14430 12804
rect 14461 12801 14473 12804
rect 14507 12801 14519 12835
rect 14461 12795 14519 12801
rect 14921 12835 14979 12841
rect 14921 12801 14933 12835
rect 14967 12832 14979 12835
rect 14967 12804 15424 12832
rect 14967 12801 14979 12804
rect 14921 12795 14979 12801
rect 14001 12767 14059 12773
rect 14001 12764 14013 12767
rect 13740 12736 14013 12764
rect 14001 12733 14013 12736
rect 14047 12733 14059 12767
rect 14001 12727 14059 12733
rect 13081 12699 13139 12705
rect 13081 12696 13093 12699
rect 12636 12668 13093 12696
rect 13081 12665 13093 12668
rect 13127 12665 13139 12699
rect 15105 12699 15163 12705
rect 15105 12696 15117 12699
rect 13081 12659 13139 12665
rect 13188 12668 15117 12696
rect 3142 12588 3148 12640
rect 3200 12628 3206 12640
rect 6641 12631 6699 12637
rect 6641 12628 6653 12631
rect 3200 12600 6653 12628
rect 3200 12588 3206 12600
rect 6641 12597 6653 12600
rect 6687 12597 6699 12631
rect 6641 12591 6699 12597
rect 11238 12588 11244 12640
rect 11296 12628 11302 12640
rect 13188 12628 13216 12668
rect 15105 12665 15117 12668
rect 15151 12665 15163 12699
rect 15396 12696 15424 12804
rect 15562 12792 15568 12844
rect 15620 12792 15626 12844
rect 15746 12792 15752 12844
rect 15804 12832 15810 12844
rect 16114 12832 16120 12844
rect 15804 12804 16120 12832
rect 15804 12792 15810 12804
rect 16114 12792 16120 12804
rect 16172 12792 16178 12844
rect 16390 12792 16396 12844
rect 16448 12792 16454 12844
rect 16758 12792 16764 12844
rect 16816 12832 16822 12844
rect 16853 12835 16911 12841
rect 16853 12832 16865 12835
rect 16816 12804 16865 12832
rect 16816 12792 16822 12804
rect 16853 12801 16865 12804
rect 16899 12801 16911 12835
rect 16853 12795 16911 12801
rect 16942 12792 16948 12844
rect 17000 12792 17006 12844
rect 15473 12767 15531 12773
rect 15473 12733 15485 12767
rect 15519 12764 15531 12767
rect 15654 12764 15660 12776
rect 15519 12736 15660 12764
rect 15519 12733 15531 12736
rect 15473 12727 15531 12733
rect 15654 12724 15660 12736
rect 15712 12724 15718 12776
rect 16574 12724 16580 12776
rect 16632 12764 16638 12776
rect 17313 12767 17371 12773
rect 17313 12764 17325 12767
rect 16632 12736 17325 12764
rect 16632 12724 16638 12736
rect 17313 12733 17325 12736
rect 17359 12733 17371 12767
rect 17313 12727 17371 12733
rect 15838 12696 15844 12708
rect 15396 12668 15844 12696
rect 15105 12659 15163 12665
rect 15838 12656 15844 12668
rect 15896 12656 15902 12708
rect 11296 12600 13216 12628
rect 11296 12588 11302 12600
rect 13906 12588 13912 12640
rect 13964 12628 13970 12640
rect 15381 12631 15439 12637
rect 15381 12628 15393 12631
rect 13964 12600 15393 12628
rect 13964 12588 13970 12600
rect 15381 12597 15393 12600
rect 15427 12628 15439 12631
rect 16206 12628 16212 12640
rect 15427 12600 16212 12628
rect 15427 12597 15439 12600
rect 15381 12591 15439 12597
rect 16206 12588 16212 12600
rect 16264 12628 16270 12640
rect 16669 12631 16727 12637
rect 16669 12628 16681 12631
rect 16264 12600 16681 12628
rect 16264 12588 16270 12600
rect 16669 12597 16681 12600
rect 16715 12597 16727 12631
rect 16669 12591 16727 12597
rect 1104 12538 17848 12560
rect 1104 12486 1918 12538
rect 1970 12486 1982 12538
rect 2034 12486 2046 12538
rect 2098 12486 2110 12538
rect 2162 12486 2174 12538
rect 2226 12486 2238 12538
rect 2290 12486 7918 12538
rect 7970 12486 7982 12538
rect 8034 12486 8046 12538
rect 8098 12486 8110 12538
rect 8162 12486 8174 12538
rect 8226 12486 8238 12538
rect 8290 12486 13918 12538
rect 13970 12486 13982 12538
rect 14034 12486 14046 12538
rect 14098 12486 14110 12538
rect 14162 12486 14174 12538
rect 14226 12486 14238 12538
rect 14290 12486 17848 12538
rect 1104 12464 17848 12486
rect 2225 12427 2283 12433
rect 2225 12393 2237 12427
rect 2271 12424 2283 12427
rect 2314 12424 2320 12436
rect 2271 12396 2320 12424
rect 2271 12393 2283 12396
rect 2225 12387 2283 12393
rect 2314 12384 2320 12396
rect 2372 12384 2378 12436
rect 3145 12427 3203 12433
rect 3145 12393 3157 12427
rect 3191 12424 3203 12427
rect 3418 12424 3424 12436
rect 3191 12396 3424 12424
rect 3191 12393 3203 12396
rect 3145 12387 3203 12393
rect 3418 12384 3424 12396
rect 3476 12384 3482 12436
rect 4062 12384 4068 12436
rect 4120 12384 4126 12436
rect 4706 12384 4712 12436
rect 4764 12384 4770 12436
rect 5626 12384 5632 12436
rect 5684 12424 5690 12436
rect 5905 12427 5963 12433
rect 5905 12424 5917 12427
rect 5684 12396 5917 12424
rect 5684 12384 5690 12396
rect 5905 12393 5917 12396
rect 5951 12393 5963 12427
rect 5905 12387 5963 12393
rect 7098 12384 7104 12436
rect 7156 12384 7162 12436
rect 15562 12384 15568 12436
rect 15620 12424 15626 12436
rect 15746 12424 15752 12436
rect 15620 12396 15752 12424
rect 15620 12384 15626 12396
rect 15746 12384 15752 12396
rect 15804 12424 15810 12436
rect 16393 12427 16451 12433
rect 16393 12424 16405 12427
rect 15804 12396 16405 12424
rect 15804 12384 15810 12396
rect 16393 12393 16405 12396
rect 16439 12393 16451 12427
rect 16393 12387 16451 12393
rect 4246 12316 4252 12368
rect 4304 12316 4310 12368
rect 4724 12356 4752 12384
rect 5166 12356 5172 12368
rect 4724 12328 5172 12356
rect 5166 12316 5172 12328
rect 5224 12356 5230 12368
rect 6273 12359 6331 12365
rect 6273 12356 6285 12359
rect 5224 12328 6285 12356
rect 5224 12316 5230 12328
rect 6273 12325 6285 12328
rect 6319 12325 6331 12359
rect 7285 12359 7343 12365
rect 7285 12356 7297 12359
rect 6273 12319 6331 12325
rect 6932 12328 7297 12356
rect 4264 12288 4292 12316
rect 3344 12260 4292 12288
rect 4709 12291 4767 12297
rect 1394 12180 1400 12232
rect 1452 12220 1458 12232
rect 1581 12223 1639 12229
rect 1581 12220 1593 12223
rect 1452 12192 1593 12220
rect 1452 12180 1458 12192
rect 1581 12189 1593 12192
rect 1627 12189 1639 12223
rect 1581 12183 1639 12189
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12220 2191 12223
rect 2498 12220 2504 12232
rect 2179 12192 2504 12220
rect 2179 12189 2191 12192
rect 2133 12183 2191 12189
rect 2498 12180 2504 12192
rect 2556 12180 2562 12232
rect 3344 12229 3372 12260
rect 4709 12257 4721 12291
rect 4755 12288 4767 12291
rect 4982 12288 4988 12300
rect 4755 12260 4988 12288
rect 4755 12257 4767 12260
rect 4709 12251 4767 12257
rect 4982 12248 4988 12260
rect 5040 12248 5046 12300
rect 6932 12297 6960 12328
rect 7285 12325 7297 12328
rect 7331 12356 7343 12359
rect 7650 12356 7656 12368
rect 7331 12328 7656 12356
rect 7331 12325 7343 12328
rect 7285 12319 7343 12325
rect 7650 12316 7656 12328
rect 7708 12316 7714 12368
rect 6917 12291 6975 12297
rect 6917 12257 6929 12291
rect 6963 12257 6975 12291
rect 6917 12251 6975 12257
rect 14458 12248 14464 12300
rect 14516 12288 14522 12300
rect 16206 12288 16212 12300
rect 14516 12260 16212 12288
rect 14516 12248 14522 12260
rect 16206 12248 16212 12260
rect 16264 12288 16270 12300
rect 16942 12288 16948 12300
rect 16264 12260 16948 12288
rect 16264 12248 16270 12260
rect 3329 12223 3387 12229
rect 3329 12189 3341 12223
rect 3375 12189 3387 12223
rect 3329 12183 3387 12189
rect 3605 12223 3663 12229
rect 3605 12189 3617 12223
rect 3651 12220 3663 12223
rect 4154 12220 4160 12232
rect 3651 12192 4160 12220
rect 3651 12189 3663 12192
rect 3605 12183 3663 12189
rect 4154 12180 4160 12192
rect 4212 12180 4218 12232
rect 4249 12223 4307 12229
rect 4249 12189 4261 12223
rect 4295 12189 4307 12223
rect 4249 12183 4307 12189
rect 4341 12223 4399 12229
rect 4341 12189 4353 12223
rect 4387 12220 4399 12223
rect 4522 12220 4528 12232
rect 4387 12192 4528 12220
rect 4387 12189 4399 12192
rect 4341 12183 4399 12189
rect 3694 12112 3700 12164
rect 3752 12152 3758 12164
rect 4264 12152 4292 12183
rect 4522 12180 4528 12192
rect 4580 12180 4586 12232
rect 5905 12223 5963 12229
rect 5905 12189 5917 12223
rect 5951 12189 5963 12223
rect 5905 12183 5963 12189
rect 6089 12223 6147 12229
rect 6089 12189 6101 12223
rect 6135 12220 6147 12223
rect 6178 12220 6184 12232
rect 6135 12192 6184 12220
rect 6135 12189 6147 12192
rect 6089 12183 6147 12189
rect 3752 12124 4292 12152
rect 5920 12152 5948 12183
rect 6178 12180 6184 12192
rect 6236 12180 6242 12232
rect 16592 12229 16620 12260
rect 16942 12248 16948 12260
rect 17000 12288 17006 12300
rect 17037 12291 17095 12297
rect 17037 12288 17049 12291
rect 17000 12260 17049 12288
rect 17000 12248 17006 12260
rect 17037 12257 17049 12260
rect 17083 12257 17095 12291
rect 17037 12251 17095 12257
rect 6365 12223 6423 12229
rect 6365 12189 6377 12223
rect 6411 12220 6423 12223
rect 6825 12223 6883 12229
rect 6411 12192 6500 12220
rect 6411 12189 6423 12192
rect 6365 12183 6423 12189
rect 6472 12152 6500 12192
rect 6825 12189 6837 12223
rect 6871 12189 6883 12223
rect 6825 12183 6883 12189
rect 16393 12223 16451 12229
rect 16393 12189 16405 12223
rect 16439 12189 16451 12223
rect 16393 12183 16451 12189
rect 16577 12223 16635 12229
rect 16577 12189 16589 12223
rect 16623 12189 16635 12223
rect 16577 12183 16635 12189
rect 5920 12124 6500 12152
rect 6840 12152 6868 12183
rect 7558 12152 7564 12164
rect 6840 12124 7564 12152
rect 3752 12112 3758 12124
rect 842 12044 848 12096
rect 900 12084 906 12096
rect 1397 12087 1455 12093
rect 1397 12084 1409 12087
rect 900 12056 1409 12084
rect 900 12044 906 12056
rect 1397 12053 1409 12056
rect 1443 12053 1455 12087
rect 1397 12047 1455 12053
rect 3513 12087 3571 12093
rect 3513 12053 3525 12087
rect 3559 12084 3571 12087
rect 4338 12084 4344 12096
rect 3559 12056 4344 12084
rect 3559 12053 3571 12056
rect 3513 12047 3571 12053
rect 4338 12044 4344 12056
rect 4396 12044 4402 12096
rect 6472 12093 6500 12124
rect 7558 12112 7564 12124
rect 7616 12112 7622 12164
rect 16408 12152 16436 12183
rect 16758 12180 16764 12232
rect 16816 12220 16822 12232
rect 16853 12223 16911 12229
rect 16853 12220 16865 12223
rect 16816 12192 16865 12220
rect 16816 12180 16822 12192
rect 16853 12189 16865 12192
rect 16899 12189 16911 12223
rect 16853 12183 16911 12189
rect 16776 12152 16804 12180
rect 16408 12124 16804 12152
rect 6457 12087 6515 12093
rect 6457 12053 6469 12087
rect 6503 12053 6515 12087
rect 6457 12047 6515 12053
rect 6638 12044 6644 12096
rect 6696 12084 6702 12096
rect 12526 12084 12532 12096
rect 6696 12056 12532 12084
rect 6696 12044 6702 12056
rect 12526 12044 12532 12056
rect 12584 12084 12590 12096
rect 13170 12084 13176 12096
rect 12584 12056 13176 12084
rect 12584 12044 12590 12056
rect 13170 12044 13176 12056
rect 13228 12044 13234 12096
rect 15654 12044 15660 12096
rect 15712 12084 15718 12096
rect 16114 12084 16120 12096
rect 15712 12056 16120 12084
rect 15712 12044 15718 12056
rect 16114 12044 16120 12056
rect 16172 12084 16178 12096
rect 16669 12087 16727 12093
rect 16669 12084 16681 12087
rect 16172 12056 16681 12084
rect 16172 12044 16178 12056
rect 16669 12053 16681 12056
rect 16715 12053 16727 12087
rect 16669 12047 16727 12053
rect 1104 11994 17848 12016
rect 1104 11942 2658 11994
rect 2710 11942 2722 11994
rect 2774 11942 2786 11994
rect 2838 11942 2850 11994
rect 2902 11942 2914 11994
rect 2966 11942 2978 11994
rect 3030 11942 8658 11994
rect 8710 11942 8722 11994
rect 8774 11942 8786 11994
rect 8838 11942 8850 11994
rect 8902 11942 8914 11994
rect 8966 11942 8978 11994
rect 9030 11942 14658 11994
rect 14710 11942 14722 11994
rect 14774 11942 14786 11994
rect 14838 11942 14850 11994
rect 14902 11942 14914 11994
rect 14966 11942 14978 11994
rect 15030 11942 17848 11994
rect 1104 11920 17848 11942
rect 3602 11840 3608 11892
rect 3660 11840 3666 11892
rect 3697 11883 3755 11889
rect 3697 11849 3709 11883
rect 3743 11880 3755 11883
rect 4338 11880 4344 11892
rect 3743 11852 4344 11880
rect 3743 11849 3755 11852
rect 3697 11843 3755 11849
rect 4338 11840 4344 11852
rect 4396 11880 4402 11892
rect 5442 11880 5448 11892
rect 4396 11852 5448 11880
rect 4396 11840 4402 11852
rect 5442 11840 5448 11852
rect 5500 11840 5506 11892
rect 6178 11840 6184 11892
rect 6236 11880 6242 11892
rect 7009 11883 7067 11889
rect 7009 11880 7021 11883
rect 6236 11852 7021 11880
rect 6236 11840 6242 11852
rect 7009 11849 7021 11852
rect 7055 11849 7067 11883
rect 7009 11843 7067 11849
rect 7558 11840 7564 11892
rect 7616 11880 7622 11892
rect 8021 11883 8079 11889
rect 8021 11880 8033 11883
rect 7616 11852 8033 11880
rect 7616 11840 7622 11852
rect 8021 11849 8033 11852
rect 8067 11849 8079 11883
rect 10781 11883 10839 11889
rect 10781 11880 10793 11883
rect 8021 11843 8079 11849
rect 9140 11852 10793 11880
rect 4433 11815 4491 11821
rect 4433 11812 4445 11815
rect 4172 11784 4445 11812
rect 4172 11756 4200 11784
rect 4433 11781 4445 11784
rect 4479 11781 4491 11815
rect 4709 11815 4767 11821
rect 4709 11812 4721 11815
rect 4433 11775 4491 11781
rect 4540 11784 4721 11812
rect 4540 11756 4568 11784
rect 4709 11781 4721 11784
rect 4755 11781 4767 11815
rect 8573 11815 8631 11821
rect 8573 11812 8585 11815
rect 4709 11775 4767 11781
rect 8220 11784 8585 11812
rect 3329 11747 3387 11753
rect 3329 11713 3341 11747
rect 3375 11744 3387 11747
rect 3418 11744 3424 11756
rect 3375 11716 3424 11744
rect 3375 11713 3387 11716
rect 3329 11707 3387 11713
rect 3418 11704 3424 11716
rect 3476 11704 3482 11756
rect 3789 11747 3847 11753
rect 3789 11713 3801 11747
rect 3835 11744 3847 11747
rect 3881 11747 3939 11753
rect 3881 11744 3893 11747
rect 3835 11716 3893 11744
rect 3835 11713 3847 11716
rect 3789 11707 3847 11713
rect 3881 11713 3893 11716
rect 3927 11713 3939 11747
rect 3881 11707 3939 11713
rect 4065 11747 4123 11753
rect 4065 11713 4077 11747
rect 4111 11713 4123 11747
rect 4065 11707 4123 11713
rect 4080 11676 4108 11707
rect 4154 11704 4160 11756
rect 4212 11704 4218 11756
rect 4341 11747 4399 11753
rect 4341 11713 4353 11747
rect 4387 11713 4399 11747
rect 4341 11707 4399 11713
rect 4246 11676 4252 11688
rect 4080 11648 4252 11676
rect 4246 11636 4252 11648
rect 4304 11636 4310 11688
rect 3694 11568 3700 11620
rect 3752 11608 3758 11620
rect 4356 11608 4384 11707
rect 4522 11704 4528 11756
rect 4580 11704 4586 11756
rect 4617 11747 4675 11753
rect 4617 11713 4629 11747
rect 4663 11744 4675 11747
rect 4798 11744 4804 11756
rect 4663 11716 4804 11744
rect 4663 11713 4675 11716
rect 4617 11707 4675 11713
rect 4798 11704 4804 11716
rect 4856 11704 4862 11756
rect 6914 11704 6920 11756
rect 6972 11704 6978 11756
rect 7006 11704 7012 11756
rect 7064 11744 7070 11756
rect 8220 11753 8248 11784
rect 8573 11781 8585 11784
rect 8619 11781 8631 11815
rect 9140 11812 9168 11852
rect 10781 11849 10793 11852
rect 10827 11849 10839 11883
rect 10781 11843 10839 11849
rect 12710 11840 12716 11892
rect 12768 11880 12774 11892
rect 13078 11880 13084 11892
rect 12768 11852 13084 11880
rect 12768 11840 12774 11852
rect 13078 11840 13084 11852
rect 13136 11880 13142 11892
rect 14369 11883 14427 11889
rect 13136 11852 13308 11880
rect 13136 11840 13142 11852
rect 8573 11775 8631 11781
rect 8680 11784 9168 11812
rect 7101 11747 7159 11753
rect 7101 11744 7113 11747
rect 7064 11716 7113 11744
rect 7064 11704 7070 11716
rect 7101 11713 7113 11716
rect 7147 11713 7159 11747
rect 7101 11707 7159 11713
rect 8205 11747 8263 11753
rect 8205 11713 8217 11747
rect 8251 11713 8263 11747
rect 8205 11707 8263 11713
rect 8386 11704 8392 11756
rect 8444 11704 8450 11756
rect 8478 11704 8484 11756
rect 8536 11744 8542 11756
rect 8680 11744 8708 11784
rect 8536 11716 8708 11744
rect 8757 11747 8815 11753
rect 8536 11704 8542 11716
rect 8757 11713 8769 11747
rect 8803 11744 8815 11747
rect 8846 11744 8852 11756
rect 8803 11716 8852 11744
rect 8803 11713 8815 11716
rect 8757 11707 8815 11713
rect 8846 11704 8852 11716
rect 8904 11704 8910 11756
rect 9033 11747 9091 11753
rect 9033 11713 9045 11747
rect 9079 11744 9091 11747
rect 9140 11744 9168 11784
rect 10137 11815 10195 11821
rect 10137 11781 10149 11815
rect 10183 11812 10195 11815
rect 11517 11815 11575 11821
rect 11517 11812 11529 11815
rect 10183 11784 11529 11812
rect 10183 11781 10195 11784
rect 10137 11775 10195 11781
rect 11517 11781 11529 11784
rect 11563 11781 11575 11815
rect 11517 11775 11575 11781
rect 11606 11772 11612 11824
rect 11664 11812 11670 11824
rect 13173 11815 13231 11821
rect 13173 11812 13185 11815
rect 11664 11784 12020 11812
rect 11664 11772 11670 11784
rect 9079 11716 9168 11744
rect 9217 11747 9275 11753
rect 9079 11713 9091 11716
rect 9033 11707 9091 11713
rect 9217 11713 9229 11747
rect 9263 11744 9275 11747
rect 9766 11744 9772 11756
rect 9263 11716 9772 11744
rect 9263 11713 9275 11716
rect 9217 11707 9275 11713
rect 3752 11580 4384 11608
rect 3752 11568 3758 11580
rect 8386 11568 8392 11620
rect 8444 11608 8450 11620
rect 9232 11608 9260 11707
rect 9766 11704 9772 11716
rect 9824 11704 9830 11756
rect 10321 11747 10379 11753
rect 10321 11713 10333 11747
rect 10367 11713 10379 11747
rect 10321 11707 10379 11713
rect 10413 11747 10471 11753
rect 10413 11713 10425 11747
rect 10459 11744 10471 11747
rect 10502 11744 10508 11756
rect 10459 11716 10508 11744
rect 10459 11713 10471 11716
rect 10413 11707 10471 11713
rect 8444 11580 9260 11608
rect 8444 11568 8450 11580
rect 9306 11568 9312 11620
rect 9364 11608 9370 11620
rect 10137 11611 10195 11617
rect 10137 11608 10149 11611
rect 9364 11580 10149 11608
rect 9364 11568 9370 11580
rect 10137 11577 10149 11580
rect 10183 11577 10195 11611
rect 10336 11608 10364 11707
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 10778 11704 10784 11756
rect 10836 11744 10842 11756
rect 11992 11753 12020 11784
rect 13004 11784 13185 11812
rect 11149 11747 11207 11753
rect 11149 11744 11161 11747
rect 10836 11716 11161 11744
rect 10836 11704 10842 11716
rect 11149 11713 11161 11716
rect 11195 11713 11207 11747
rect 11149 11707 11207 11713
rect 11701 11747 11759 11753
rect 11701 11713 11713 11747
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 11977 11747 12035 11753
rect 11977 11713 11989 11747
rect 12023 11713 12035 11747
rect 11977 11707 12035 11713
rect 12437 11747 12495 11753
rect 12437 11713 12449 11747
rect 12483 11744 12495 11747
rect 12526 11744 12532 11756
rect 12483 11716 12532 11744
rect 12483 11713 12495 11716
rect 12437 11707 12495 11713
rect 11241 11679 11299 11685
rect 11241 11645 11253 11679
rect 11287 11676 11299 11679
rect 11716 11676 11744 11707
rect 12526 11704 12532 11716
rect 12584 11704 12590 11756
rect 12710 11704 12716 11756
rect 12768 11704 12774 11756
rect 12805 11747 12863 11753
rect 12805 11713 12817 11747
rect 12851 11744 12863 11747
rect 12894 11744 12900 11756
rect 12851 11716 12900 11744
rect 12851 11713 12863 11716
rect 12805 11707 12863 11713
rect 12894 11704 12900 11716
rect 12952 11704 12958 11756
rect 13004 11753 13032 11784
rect 13173 11781 13185 11784
rect 13219 11781 13231 11815
rect 13173 11775 13231 11781
rect 13280 11753 13308 11852
rect 14369 11849 14381 11883
rect 14415 11880 14427 11883
rect 14645 11883 14703 11889
rect 14645 11880 14657 11883
rect 14415 11852 14657 11880
rect 14415 11849 14427 11852
rect 14369 11843 14427 11849
rect 14645 11849 14657 11852
rect 14691 11849 14703 11883
rect 14645 11843 14703 11849
rect 15488 11852 15792 11880
rect 13909 11815 13967 11821
rect 13909 11781 13921 11815
rect 13955 11812 13967 11815
rect 15286 11812 15292 11824
rect 13955 11784 15292 11812
rect 13955 11781 13967 11784
rect 13909 11775 13967 11781
rect 15286 11772 15292 11784
rect 15344 11772 15350 11824
rect 12989 11747 13047 11753
rect 12989 11713 13001 11747
rect 13035 11713 13047 11747
rect 12989 11707 13047 11713
rect 13081 11747 13139 11753
rect 13081 11713 13093 11747
rect 13127 11713 13139 11747
rect 13081 11707 13139 11713
rect 13265 11747 13323 11753
rect 13265 11713 13277 11747
rect 13311 11713 13323 11747
rect 13265 11707 13323 11713
rect 14001 11747 14059 11753
rect 14001 11713 14013 11747
rect 14047 11744 14059 11747
rect 14550 11744 14556 11756
rect 14047 11716 14556 11744
rect 14047 11713 14059 11716
rect 14001 11707 14059 11713
rect 11287 11648 11744 11676
rect 11287 11645 11299 11648
rect 11241 11639 11299 11645
rect 11606 11608 11612 11620
rect 10336 11580 11612 11608
rect 10137 11571 10195 11577
rect 11606 11568 11612 11580
rect 11664 11568 11670 11620
rect 11716 11608 11744 11648
rect 12618 11636 12624 11688
rect 12676 11636 12682 11688
rect 13096 11676 13124 11707
rect 14550 11704 14556 11716
rect 14608 11704 14614 11756
rect 15488 11753 15516 11852
rect 15764 11812 15792 11852
rect 15838 11840 15844 11892
rect 15896 11880 15902 11892
rect 16117 11883 16175 11889
rect 16117 11880 16129 11883
rect 15896 11852 16129 11880
rect 15896 11840 15902 11852
rect 16117 11849 16129 11852
rect 16163 11849 16175 11883
rect 16117 11843 16175 11849
rect 16942 11840 16948 11892
rect 17000 11840 17006 11892
rect 16574 11812 16580 11824
rect 15764 11784 16580 11812
rect 16574 11772 16580 11784
rect 16632 11812 16638 11824
rect 16960 11812 16988 11840
rect 16632 11784 16896 11812
rect 16960 11784 17356 11812
rect 16632 11772 16638 11784
rect 14642 11747 14700 11753
rect 14642 11713 14654 11747
rect 14688 11744 14700 11747
rect 15197 11747 15255 11753
rect 15197 11744 15209 11747
rect 14688 11716 15209 11744
rect 14688 11713 14700 11716
rect 14642 11707 14700 11713
rect 15197 11713 15209 11716
rect 15243 11713 15255 11747
rect 15197 11707 15255 11713
rect 15381 11747 15439 11753
rect 15381 11713 15393 11747
rect 15427 11713 15439 11747
rect 15381 11707 15439 11713
rect 15473 11747 15531 11753
rect 15473 11713 15485 11747
rect 15519 11713 15531 11747
rect 15473 11707 15531 11713
rect 13170 11676 13176 11688
rect 13096 11648 13176 11676
rect 13170 11636 13176 11648
rect 13228 11636 13234 11688
rect 13446 11636 13452 11688
rect 13504 11676 13510 11688
rect 13725 11679 13783 11685
rect 13725 11676 13737 11679
rect 13504 11648 13737 11676
rect 13504 11636 13510 11648
rect 13725 11645 13737 11648
rect 13771 11645 13783 11679
rect 13725 11639 13783 11645
rect 15102 11636 15108 11688
rect 15160 11636 15166 11688
rect 15396 11676 15424 11707
rect 15654 11704 15660 11756
rect 15712 11704 15718 11756
rect 15746 11704 15752 11756
rect 15804 11704 15810 11756
rect 15841 11747 15899 11753
rect 15841 11713 15853 11747
rect 15887 11744 15899 11747
rect 16022 11744 16028 11756
rect 15887 11716 16028 11744
rect 15887 11713 15899 11716
rect 15841 11707 15899 11713
rect 15856 11676 15884 11707
rect 16022 11704 16028 11716
rect 16080 11704 16086 11756
rect 16206 11704 16212 11756
rect 16264 11744 16270 11756
rect 16301 11747 16359 11753
rect 16301 11744 16313 11747
rect 16264 11716 16313 11744
rect 16264 11704 16270 11716
rect 16301 11713 16313 11716
rect 16347 11713 16359 11747
rect 16301 11707 16359 11713
rect 16485 11747 16543 11753
rect 16485 11713 16497 11747
rect 16531 11744 16543 11747
rect 16758 11744 16764 11756
rect 16531 11716 16764 11744
rect 16531 11713 16543 11716
rect 16485 11707 16543 11713
rect 16758 11704 16764 11716
rect 16816 11704 16822 11756
rect 16868 11753 16896 11784
rect 16853 11747 16911 11753
rect 16853 11713 16865 11747
rect 16899 11744 16911 11747
rect 16942 11744 16948 11756
rect 16899 11716 16948 11744
rect 16899 11713 16911 11716
rect 16853 11707 16911 11713
rect 16942 11704 16948 11716
rect 17000 11704 17006 11756
rect 17328 11753 17356 11784
rect 17129 11747 17187 11753
rect 17129 11713 17141 11747
rect 17175 11713 17187 11747
rect 17129 11707 17187 11713
rect 17313 11747 17371 11753
rect 17313 11713 17325 11747
rect 17359 11713 17371 11747
rect 17313 11707 17371 11713
rect 15396 11648 15884 11676
rect 16117 11679 16175 11685
rect 14461 11611 14519 11617
rect 14461 11608 14473 11611
rect 11716 11580 14473 11608
rect 14461 11577 14473 11580
rect 14507 11577 14519 11611
rect 15396 11608 15424 11648
rect 16117 11645 16129 11679
rect 16163 11676 16175 11679
rect 16776 11676 16804 11704
rect 17144 11676 17172 11707
rect 16163 11648 16712 11676
rect 16776 11648 17172 11676
rect 16163 11645 16175 11648
rect 16117 11639 16175 11645
rect 14461 11571 14519 11577
rect 15028 11580 15424 11608
rect 11698 11500 11704 11552
rect 11756 11540 11762 11552
rect 11885 11543 11943 11549
rect 11885 11540 11897 11543
rect 11756 11512 11897 11540
rect 11756 11500 11762 11512
rect 11885 11509 11897 11512
rect 11931 11509 11943 11543
rect 11885 11503 11943 11509
rect 12253 11543 12311 11549
rect 12253 11509 12265 11543
rect 12299 11540 12311 11543
rect 12986 11540 12992 11552
rect 12299 11512 12992 11540
rect 12299 11509 12311 11512
rect 12253 11503 12311 11509
rect 12986 11500 12992 11512
rect 13044 11500 13050 11552
rect 13630 11500 13636 11552
rect 13688 11540 13694 11552
rect 15028 11549 15056 11580
rect 15013 11543 15071 11549
rect 15013 11540 15025 11543
rect 13688 11512 15025 11540
rect 13688 11500 13694 11512
rect 15013 11509 15025 11512
rect 15059 11509 15071 11543
rect 15013 11503 15071 11509
rect 15654 11500 15660 11552
rect 15712 11540 15718 11552
rect 16684 11549 16712 11648
rect 15933 11543 15991 11549
rect 15933 11540 15945 11543
rect 15712 11512 15945 11540
rect 15712 11500 15718 11512
rect 15933 11509 15945 11512
rect 15979 11540 15991 11543
rect 16393 11543 16451 11549
rect 16393 11540 16405 11543
rect 15979 11512 16405 11540
rect 15979 11509 15991 11512
rect 15933 11503 15991 11509
rect 16393 11509 16405 11512
rect 16439 11509 16451 11543
rect 16393 11503 16451 11509
rect 16669 11543 16727 11549
rect 16669 11509 16681 11543
rect 16715 11540 16727 11543
rect 17034 11540 17040 11552
rect 16715 11512 17040 11540
rect 16715 11509 16727 11512
rect 16669 11503 16727 11509
rect 17034 11500 17040 11512
rect 17092 11500 17098 11552
rect 1104 11450 17848 11472
rect 1104 11398 1918 11450
rect 1970 11398 1982 11450
rect 2034 11398 2046 11450
rect 2098 11398 2110 11450
rect 2162 11398 2174 11450
rect 2226 11398 2238 11450
rect 2290 11398 7918 11450
rect 7970 11398 7982 11450
rect 8034 11398 8046 11450
rect 8098 11398 8110 11450
rect 8162 11398 8174 11450
rect 8226 11398 8238 11450
rect 8290 11398 13918 11450
rect 13970 11398 13982 11450
rect 14034 11398 14046 11450
rect 14098 11398 14110 11450
rect 14162 11398 14174 11450
rect 14226 11398 14238 11450
rect 14290 11398 17848 11450
rect 1104 11376 17848 11398
rect 1394 11296 1400 11348
rect 1452 11296 1458 11348
rect 4798 11296 4804 11348
rect 4856 11296 4862 11348
rect 5442 11296 5448 11348
rect 5500 11296 5506 11348
rect 10778 11296 10784 11348
rect 10836 11296 10842 11348
rect 15654 11296 15660 11348
rect 15712 11296 15718 11348
rect 3789 11271 3847 11277
rect 3789 11268 3801 11271
rect 3068 11240 3801 11268
rect 2869 11203 2927 11209
rect 2869 11169 2881 11203
rect 2915 11200 2927 11203
rect 3068 11200 3096 11240
rect 3789 11237 3801 11240
rect 3835 11237 3847 11271
rect 3789 11231 3847 11237
rect 2915 11172 3096 11200
rect 2915 11169 2927 11172
rect 2869 11163 2927 11169
rect 3142 11160 3148 11212
rect 3200 11160 3206 11212
rect 3694 11160 3700 11212
rect 3752 11200 3758 11212
rect 4249 11203 4307 11209
rect 4249 11200 4261 11203
rect 3752 11172 4261 11200
rect 3752 11160 3758 11172
rect 4249 11169 4261 11172
rect 4295 11169 4307 11203
rect 4249 11163 4307 11169
rect 3421 11135 3479 11141
rect 3421 11101 3433 11135
rect 3467 11101 3479 11135
rect 3421 11095 3479 11101
rect 4157 11135 4215 11141
rect 4157 11101 4169 11135
rect 4203 11132 4215 11135
rect 4816 11132 4844 11296
rect 6914 11228 6920 11280
rect 6972 11268 6978 11280
rect 8941 11271 8999 11277
rect 8941 11268 8953 11271
rect 6972 11240 8953 11268
rect 6972 11228 6978 11240
rect 7116 11209 7144 11240
rect 8941 11237 8953 11240
rect 8987 11237 8999 11271
rect 16114 11268 16120 11280
rect 8941 11231 8999 11237
rect 12728 11240 14504 11268
rect 12728 11212 12756 11240
rect 5169 11203 5227 11209
rect 5169 11169 5181 11203
rect 5215 11200 5227 11203
rect 6641 11203 6699 11209
rect 5215 11172 5580 11200
rect 5215 11169 5227 11172
rect 5169 11163 5227 11169
rect 5552 11141 5580 11172
rect 6641 11169 6653 11203
rect 6687 11169 6699 11203
rect 6641 11163 6699 11169
rect 7101 11203 7159 11209
rect 7101 11169 7113 11203
rect 7147 11169 7159 11203
rect 7101 11163 7159 11169
rect 4203 11104 4844 11132
rect 5077 11135 5135 11141
rect 4203 11101 4215 11104
rect 4157 11095 4215 11101
rect 5077 11101 5089 11135
rect 5123 11132 5135 11135
rect 5353 11135 5411 11141
rect 5353 11132 5365 11135
rect 5123 11104 5365 11132
rect 5123 11101 5135 11104
rect 5077 11095 5135 11101
rect 5353 11101 5365 11104
rect 5399 11101 5411 11135
rect 5353 11095 5411 11101
rect 5537 11135 5595 11141
rect 5537 11101 5549 11135
rect 5583 11132 5595 11135
rect 6656 11132 6684 11163
rect 8478 11160 8484 11212
rect 8536 11160 8542 11212
rect 8757 11203 8815 11209
rect 8757 11169 8769 11203
rect 8803 11200 8815 11203
rect 9217 11203 9275 11209
rect 9217 11200 9229 11203
rect 8803 11172 9229 11200
rect 8803 11169 8815 11172
rect 8757 11163 8815 11169
rect 9217 11169 9229 11172
rect 9263 11169 9275 11203
rect 9217 11163 9275 11169
rect 10502 11160 10508 11212
rect 10560 11200 10566 11212
rect 11698 11200 11704 11212
rect 10560 11172 11704 11200
rect 10560 11160 10566 11172
rect 11698 11160 11704 11172
rect 11756 11160 11762 11212
rect 12621 11203 12679 11209
rect 12621 11169 12633 11203
rect 12667 11200 12679 11203
rect 12710 11200 12716 11212
rect 12667 11172 12716 11200
rect 12667 11169 12679 11172
rect 12621 11163 12679 11169
rect 12710 11160 12716 11172
rect 12768 11160 12774 11212
rect 12986 11160 12992 11212
rect 13044 11160 13050 11212
rect 13357 11203 13415 11209
rect 13357 11169 13369 11203
rect 13403 11200 13415 11203
rect 14366 11200 14372 11212
rect 13403 11172 14372 11200
rect 13403 11169 13415 11172
rect 13357 11163 13415 11169
rect 14366 11160 14372 11172
rect 14424 11160 14430 11212
rect 14476 11200 14504 11240
rect 15120 11240 16120 11268
rect 15120 11209 15148 11240
rect 16114 11228 16120 11240
rect 16172 11228 16178 11280
rect 15105 11203 15163 11209
rect 14476 11172 15056 11200
rect 5583 11104 6684 11132
rect 5583 11101 5595 11104
rect 5537 11095 5595 11101
rect 3329 11067 3387 11073
rect 3329 11064 3341 11067
rect 2438 11036 3341 11064
rect 3329 11033 3341 11036
rect 3375 11033 3387 11067
rect 3329 11027 3387 11033
rect 2498 10956 2504 11008
rect 2556 10996 2562 11008
rect 3436 10996 3464 11095
rect 5368 11064 5396 11095
rect 7006 11092 7012 11144
rect 7064 11092 7070 11144
rect 8386 11092 8392 11144
rect 8444 11092 8450 11144
rect 8846 11092 8852 11144
rect 8904 11132 8910 11144
rect 9309 11135 9367 11141
rect 9309 11132 9321 11135
rect 8904 11104 9321 11132
rect 8904 11092 8910 11104
rect 9309 11101 9321 11104
rect 9355 11101 9367 11135
rect 9309 11095 9367 11101
rect 10413 11135 10471 11141
rect 10413 11101 10425 11135
rect 10459 11132 10471 11135
rect 11606 11132 11612 11144
rect 10459 11104 11612 11132
rect 10459 11101 10471 11104
rect 10413 11095 10471 11101
rect 6914 11064 6920 11076
rect 5368 11036 6920 11064
rect 6914 11024 6920 11036
rect 6972 11024 6978 11076
rect 7024 11064 7052 11092
rect 8478 11064 8484 11076
rect 7024 11036 8484 11064
rect 8478 11024 8484 11036
rect 8536 11024 8542 11076
rect 9324 11064 9352 11095
rect 11606 11092 11612 11104
rect 11664 11092 11670 11144
rect 12434 11092 12440 11144
rect 12492 11132 12498 11144
rect 12529 11135 12587 11141
rect 12529 11132 12541 11135
rect 12492 11104 12541 11132
rect 12492 11092 12498 11104
rect 12529 11101 12541 11104
rect 12575 11132 12587 11135
rect 13262 11132 13268 11144
rect 12575 11104 13268 11132
rect 12575 11101 12587 11104
rect 12529 11095 12587 11101
rect 13262 11092 13268 11104
rect 13320 11092 13326 11144
rect 13446 11092 13452 11144
rect 13504 11132 13510 11144
rect 13541 11135 13599 11141
rect 13541 11132 13553 11135
rect 13504 11104 13553 11132
rect 13504 11092 13510 11104
rect 13541 11101 13553 11104
rect 13587 11101 13599 11135
rect 13541 11095 13599 11101
rect 13909 11135 13967 11141
rect 13909 11101 13921 11135
rect 13955 11132 13967 11135
rect 14737 11135 14795 11141
rect 14737 11132 14749 11135
rect 13955 11104 14749 11132
rect 13955 11101 13967 11104
rect 13909 11095 13967 11101
rect 14737 11101 14749 11104
rect 14783 11101 14795 11135
rect 14737 11095 14795 11101
rect 14921 11135 14979 11141
rect 14921 11101 14933 11135
rect 14967 11101 14979 11135
rect 15028 11132 15056 11172
rect 15105 11169 15117 11203
rect 15151 11169 15163 11203
rect 15378 11200 15384 11212
rect 15105 11163 15163 11169
rect 15212 11172 15384 11200
rect 15212 11141 15240 11172
rect 15378 11160 15384 11172
rect 15436 11200 15442 11212
rect 15841 11203 15899 11209
rect 15436 11172 15608 11200
rect 15436 11160 15442 11172
rect 15197 11135 15255 11141
rect 15197 11132 15209 11135
rect 15028 11104 15209 11132
rect 14921 11095 14979 11101
rect 15197 11101 15209 11104
rect 15243 11101 15255 11135
rect 15197 11095 15255 11101
rect 12345 11067 12403 11073
rect 12345 11064 12357 11067
rect 9324 11036 12357 11064
rect 12345 11033 12357 11036
rect 12391 11033 12403 11067
rect 12345 11027 12403 11033
rect 12912 11036 13124 11064
rect 2556 10968 3464 10996
rect 2556 10956 2562 10968
rect 10686 10956 10692 11008
rect 10744 10996 10750 11008
rect 12912 10996 12940 11036
rect 10744 10968 12940 10996
rect 13096 10996 13124 11036
rect 13354 11024 13360 11076
rect 13412 11064 13418 11076
rect 13722 11064 13728 11076
rect 13412 11036 13728 11064
rect 13412 11024 13418 11036
rect 13722 11024 13728 11036
rect 13780 11064 13786 11076
rect 14936 11064 14964 11095
rect 15286 11092 15292 11144
rect 15344 11092 15350 11144
rect 15580 11141 15608 11172
rect 15841 11169 15853 11203
rect 15887 11200 15899 11203
rect 17034 11200 17040 11212
rect 15887 11172 17040 11200
rect 15887 11169 15899 11172
rect 15841 11163 15899 11169
rect 17034 11160 17040 11172
rect 17092 11160 17098 11212
rect 15473 11135 15531 11141
rect 15473 11101 15485 11135
rect 15519 11101 15531 11135
rect 15473 11095 15531 11101
rect 15565 11135 15623 11141
rect 15565 11101 15577 11135
rect 15611 11101 15623 11135
rect 15565 11095 15623 11101
rect 13780 11036 14964 11064
rect 15488 11064 15516 11095
rect 15746 11092 15752 11144
rect 15804 11132 15810 11144
rect 16485 11135 16543 11141
rect 16485 11132 16497 11135
rect 15804 11104 16497 11132
rect 15804 11092 15810 11104
rect 16485 11101 16497 11104
rect 16531 11132 16543 11135
rect 16758 11132 16764 11144
rect 16531 11104 16764 11132
rect 16531 11101 16543 11104
rect 16485 11095 16543 11101
rect 16758 11092 16764 11104
rect 16816 11092 16822 11144
rect 15841 11067 15899 11073
rect 15841 11064 15853 11067
rect 15488 11036 15853 11064
rect 13780 11024 13786 11036
rect 15841 11033 15853 11036
rect 15887 11033 15899 11067
rect 15841 11027 15899 11033
rect 16114 11024 16120 11076
rect 16172 11024 16178 11076
rect 16298 11024 16304 11076
rect 16356 11024 16362 11076
rect 13541 10999 13599 11005
rect 13541 10996 13553 10999
rect 13096 10968 13553 10996
rect 10744 10956 10750 10968
rect 13541 10965 13553 10968
rect 13587 10965 13599 10999
rect 13541 10959 13599 10965
rect 1104 10906 17848 10928
rect 1104 10854 2658 10906
rect 2710 10854 2722 10906
rect 2774 10854 2786 10906
rect 2838 10854 2850 10906
rect 2902 10854 2914 10906
rect 2966 10854 2978 10906
rect 3030 10854 8658 10906
rect 8710 10854 8722 10906
rect 8774 10854 8786 10906
rect 8838 10854 8850 10906
rect 8902 10854 8914 10906
rect 8966 10854 8978 10906
rect 9030 10854 14658 10906
rect 14710 10854 14722 10906
rect 14774 10854 14786 10906
rect 14838 10854 14850 10906
rect 14902 10854 14914 10906
rect 14966 10854 14978 10906
rect 15030 10854 17848 10906
rect 1104 10832 17848 10854
rect 1302 10752 1308 10804
rect 1360 10792 1366 10804
rect 1397 10795 1455 10801
rect 1397 10792 1409 10795
rect 1360 10764 1409 10792
rect 1360 10752 1366 10764
rect 1397 10761 1409 10764
rect 1443 10761 1455 10795
rect 1397 10755 1455 10761
rect 15102 10752 15108 10804
rect 15160 10792 15166 10804
rect 15197 10795 15255 10801
rect 15197 10792 15209 10795
rect 15160 10764 15209 10792
rect 15160 10752 15166 10764
rect 15197 10761 15209 10764
rect 15243 10761 15255 10795
rect 15197 10755 15255 10761
rect 6638 10684 6644 10736
rect 6696 10724 6702 10736
rect 11241 10727 11299 10733
rect 6696 10696 7130 10724
rect 6696 10684 6702 10696
rect 11241 10693 11253 10727
rect 11287 10724 11299 10727
rect 16574 10724 16580 10736
rect 11287 10696 16580 10724
rect 11287 10693 11299 10696
rect 11241 10687 11299 10693
rect 16574 10684 16580 10696
rect 16632 10684 16638 10736
rect 1394 10616 1400 10668
rect 1452 10656 1458 10668
rect 1581 10659 1639 10665
rect 1581 10656 1593 10659
rect 1452 10628 1593 10656
rect 1452 10616 1458 10628
rect 1581 10625 1593 10628
rect 1627 10625 1639 10659
rect 1581 10619 1639 10625
rect 6362 10616 6368 10668
rect 6420 10616 6426 10668
rect 11606 10616 11612 10668
rect 11664 10656 11670 10668
rect 11701 10659 11759 10665
rect 11701 10656 11713 10659
rect 11664 10628 11713 10656
rect 11664 10616 11670 10628
rect 11701 10625 11713 10628
rect 11747 10625 11759 10659
rect 11701 10619 11759 10625
rect 11885 10659 11943 10665
rect 11885 10625 11897 10659
rect 11931 10625 11943 10659
rect 11885 10619 11943 10625
rect 15105 10659 15163 10665
rect 15105 10625 15117 10659
rect 15151 10625 15163 10659
rect 15105 10619 15163 10625
rect 15289 10659 15347 10665
rect 15289 10625 15301 10659
rect 15335 10656 15347 10659
rect 15746 10656 15752 10668
rect 15335 10628 15752 10656
rect 15335 10625 15347 10628
rect 15289 10619 15347 10625
rect 5718 10548 5724 10600
rect 5776 10588 5782 10600
rect 6641 10591 6699 10597
rect 6641 10588 6653 10591
rect 5776 10560 6653 10588
rect 5776 10548 5782 10560
rect 6641 10557 6653 10560
rect 6687 10557 6699 10591
rect 6641 10551 6699 10557
rect 7098 10548 7104 10600
rect 7156 10588 7162 10600
rect 8389 10591 8447 10597
rect 8389 10588 8401 10591
rect 7156 10560 8401 10588
rect 7156 10548 7162 10560
rect 8389 10557 8401 10560
rect 8435 10588 8447 10591
rect 10778 10588 10784 10600
rect 8435 10560 10784 10588
rect 8435 10557 8447 10560
rect 8389 10551 8447 10557
rect 10778 10548 10784 10560
rect 10836 10548 10842 10600
rect 10962 10548 10968 10600
rect 11020 10588 11026 10600
rect 11900 10588 11928 10619
rect 11020 10560 11928 10588
rect 15120 10588 15148 10619
rect 15746 10616 15752 10628
rect 15804 10656 15810 10668
rect 15804 10628 16068 10656
rect 15804 10616 15810 10628
rect 15194 10588 15200 10600
rect 15120 10560 15200 10588
rect 11020 10548 11026 10560
rect 15194 10548 15200 10560
rect 15252 10588 15258 10600
rect 15654 10588 15660 10600
rect 15252 10560 15660 10588
rect 15252 10548 15258 10560
rect 15654 10548 15660 10560
rect 15712 10548 15718 10600
rect 16040 10520 16068 10628
rect 16666 10616 16672 10668
rect 16724 10616 16730 10668
rect 16758 10616 16764 10668
rect 16816 10616 16822 10668
rect 16942 10548 16948 10600
rect 17000 10548 17006 10600
rect 17034 10520 17040 10532
rect 16040 10492 17040 10520
rect 17034 10480 17040 10492
rect 17092 10480 17098 10532
rect 9674 10412 9680 10464
rect 9732 10452 9738 10464
rect 9769 10455 9827 10461
rect 9769 10452 9781 10455
rect 9732 10424 9781 10452
rect 9732 10412 9738 10424
rect 9769 10421 9781 10424
rect 9815 10421 9827 10455
rect 9769 10415 9827 10421
rect 10870 10412 10876 10464
rect 10928 10452 10934 10464
rect 11517 10455 11575 10461
rect 11517 10452 11529 10455
rect 10928 10424 11529 10452
rect 10928 10412 10934 10424
rect 11517 10421 11529 10424
rect 11563 10421 11575 10455
rect 11517 10415 11575 10421
rect 16853 10455 16911 10461
rect 16853 10421 16865 10455
rect 16899 10452 16911 10455
rect 16942 10452 16948 10464
rect 16899 10424 16948 10452
rect 16899 10421 16911 10424
rect 16853 10415 16911 10421
rect 16942 10412 16948 10424
rect 17000 10412 17006 10464
rect 1104 10362 17848 10384
rect 1104 10310 1918 10362
rect 1970 10310 1982 10362
rect 2034 10310 2046 10362
rect 2098 10310 2110 10362
rect 2162 10310 2174 10362
rect 2226 10310 2238 10362
rect 2290 10310 7918 10362
rect 7970 10310 7982 10362
rect 8034 10310 8046 10362
rect 8098 10310 8110 10362
rect 8162 10310 8174 10362
rect 8226 10310 8238 10362
rect 8290 10310 13918 10362
rect 13970 10310 13982 10362
rect 14034 10310 14046 10362
rect 14098 10310 14110 10362
rect 14162 10310 14174 10362
rect 14226 10310 14238 10362
rect 14290 10310 17848 10362
rect 1104 10288 17848 10310
rect 1394 10208 1400 10260
rect 1452 10208 1458 10260
rect 6638 10208 6644 10260
rect 6696 10208 6702 10260
rect 12710 10208 12716 10260
rect 12768 10248 12774 10260
rect 13262 10248 13268 10260
rect 12768 10220 13268 10248
rect 12768 10208 12774 10220
rect 13262 10208 13268 10220
rect 13320 10248 13326 10260
rect 15013 10251 15071 10257
rect 13320 10220 14964 10248
rect 13320 10208 13326 10220
rect 3878 10140 3884 10192
rect 3936 10140 3942 10192
rect 9766 10140 9772 10192
rect 9824 10180 9830 10192
rect 10505 10183 10563 10189
rect 10505 10180 10517 10183
rect 9824 10152 10517 10180
rect 9824 10140 9830 10152
rect 10505 10149 10517 10152
rect 10551 10149 10563 10183
rect 10505 10143 10563 10149
rect 10778 10140 10784 10192
rect 10836 10180 10842 10192
rect 12894 10180 12900 10192
rect 10836 10152 12480 10180
rect 10836 10140 10842 10152
rect 2869 10115 2927 10121
rect 2869 10081 2881 10115
rect 2915 10112 2927 10115
rect 3789 10115 3847 10121
rect 3789 10112 3801 10115
rect 2915 10084 3801 10112
rect 2915 10081 2927 10084
rect 2869 10075 2927 10081
rect 3789 10081 3801 10084
rect 3835 10081 3847 10115
rect 3789 10075 3847 10081
rect 10229 10115 10287 10121
rect 10229 10081 10241 10115
rect 10275 10112 10287 10115
rect 10275 10084 10548 10112
rect 10275 10081 10287 10084
rect 10229 10075 10287 10081
rect 3142 10004 3148 10056
rect 3200 10004 3206 10056
rect 6549 10047 6607 10053
rect 6549 10013 6561 10047
rect 6595 10013 6607 10047
rect 6549 10007 6607 10013
rect 9953 10047 10011 10053
rect 9953 10013 9965 10047
rect 9999 10013 10011 10047
rect 9953 10007 10011 10013
rect 2406 9936 2412 9988
rect 2464 9936 2470 9988
rect 4246 9936 4252 9988
rect 4304 9936 4310 9988
rect 2498 9868 2504 9920
rect 2556 9908 2562 9920
rect 6564 9908 6592 10007
rect 9766 9936 9772 9988
rect 9824 9976 9830 9988
rect 9968 9976 9996 10007
rect 10042 10004 10048 10056
rect 10100 10004 10106 10056
rect 10520 10053 10548 10084
rect 10686 10072 10692 10124
rect 10744 10072 10750 10124
rect 10505 10047 10563 10053
rect 10505 10013 10517 10047
rect 10551 10013 10563 10047
rect 10505 10007 10563 10013
rect 10870 10004 10876 10056
rect 10928 10004 10934 10056
rect 12360 10053 12388 10152
rect 12345 10047 12403 10053
rect 12345 10013 12357 10047
rect 12391 10013 12403 10047
rect 12345 10007 12403 10013
rect 11606 9976 11612 9988
rect 9824 9948 11612 9976
rect 9824 9936 9830 9948
rect 11606 9936 11612 9948
rect 11664 9936 11670 9988
rect 12452 9976 12480 10152
rect 12544 10152 12900 10180
rect 12544 10056 12572 10152
rect 12894 10140 12900 10152
rect 12952 10140 12958 10192
rect 13630 10140 13636 10192
rect 13688 10180 13694 10192
rect 14090 10180 14096 10192
rect 13688 10152 14096 10180
rect 13688 10140 13694 10152
rect 14090 10140 14096 10152
rect 14148 10140 14154 10192
rect 14458 10140 14464 10192
rect 14516 10180 14522 10192
rect 14553 10183 14611 10189
rect 14553 10180 14565 10183
rect 14516 10152 14565 10180
rect 14516 10140 14522 10152
rect 14553 10149 14565 10152
rect 14599 10149 14611 10183
rect 14936 10180 14964 10220
rect 15013 10217 15025 10251
rect 15059 10248 15071 10251
rect 15194 10248 15200 10260
rect 15059 10220 15200 10248
rect 15059 10217 15071 10220
rect 15013 10211 15071 10217
rect 15194 10208 15200 10220
rect 15252 10208 15258 10260
rect 16393 10251 16451 10257
rect 16393 10217 16405 10251
rect 16439 10248 16451 10251
rect 16850 10248 16856 10260
rect 16439 10220 16856 10248
rect 16439 10217 16451 10220
rect 16393 10211 16451 10217
rect 16850 10208 16856 10220
rect 16908 10208 16914 10260
rect 16574 10180 16580 10192
rect 14936 10152 16580 10180
rect 14553 10143 14611 10149
rect 12636 10084 13124 10112
rect 12526 10004 12532 10056
rect 12584 10004 12590 10056
rect 12636 10053 12664 10084
rect 13096 10056 13124 10084
rect 13446 10072 13452 10124
rect 13504 10112 13510 10124
rect 15197 10115 15255 10121
rect 13504 10084 14964 10112
rect 13504 10072 13510 10084
rect 12621 10047 12679 10053
rect 12621 10013 12633 10047
rect 12667 10013 12679 10047
rect 12621 10007 12679 10013
rect 12710 10004 12716 10056
rect 12768 10044 12774 10056
rect 12805 10047 12863 10053
rect 12805 10044 12817 10047
rect 12768 10016 12817 10044
rect 12768 10004 12774 10016
rect 12805 10013 12817 10016
rect 12851 10013 12863 10047
rect 12805 10007 12863 10013
rect 12897 10047 12955 10053
rect 12897 10013 12909 10047
rect 12943 10013 12955 10047
rect 12897 10007 12955 10013
rect 12912 9976 12940 10007
rect 13078 10004 13084 10056
rect 13136 10004 13142 10056
rect 13538 10004 13544 10056
rect 13596 10044 13602 10056
rect 13906 10044 13912 10056
rect 13596 10016 13912 10044
rect 13596 10004 13602 10016
rect 13906 10004 13912 10016
rect 13964 10004 13970 10056
rect 14550 10004 14556 10056
rect 14608 10004 14614 10056
rect 14936 10053 14964 10084
rect 15197 10081 15209 10115
rect 15243 10112 15255 10115
rect 15746 10112 15752 10124
rect 15243 10084 15752 10112
rect 15243 10081 15255 10084
rect 15197 10075 15255 10081
rect 15746 10072 15752 10084
rect 15804 10072 15810 10124
rect 14829 10047 14887 10053
rect 14829 10013 14841 10047
rect 14875 10013 14887 10047
rect 14829 10007 14887 10013
rect 14921 10047 14979 10053
rect 14921 10013 14933 10047
rect 14967 10044 14979 10047
rect 15286 10044 15292 10056
rect 14967 10016 15292 10044
rect 14967 10013 14979 10016
rect 14921 10007 14979 10013
rect 12986 9976 12992 9988
rect 12452 9948 12992 9976
rect 12986 9936 12992 9948
rect 13044 9976 13050 9988
rect 13446 9976 13452 9988
rect 13044 9948 13452 9976
rect 13044 9936 13050 9948
rect 13446 9936 13452 9948
rect 13504 9936 13510 9988
rect 14844 9976 14872 10007
rect 15286 10004 15292 10016
rect 15344 10004 15350 10056
rect 15562 10004 15568 10056
rect 15620 10004 15626 10056
rect 15654 10004 15660 10056
rect 15712 10044 15718 10056
rect 16316 10053 16344 10152
rect 16574 10140 16580 10152
rect 16632 10140 16638 10192
rect 16666 10140 16672 10192
rect 16724 10140 16730 10192
rect 16209 10047 16267 10053
rect 16209 10044 16221 10047
rect 15712 10016 16221 10044
rect 15712 10004 15718 10016
rect 16209 10013 16221 10016
rect 16255 10013 16267 10047
rect 16209 10007 16267 10013
rect 16301 10047 16359 10053
rect 16301 10013 16313 10047
rect 16347 10013 16359 10047
rect 16301 10007 16359 10013
rect 16942 10004 16948 10056
rect 17000 10004 17006 10056
rect 17034 10004 17040 10056
rect 17092 10004 17098 10056
rect 17126 10004 17132 10056
rect 17184 10044 17190 10056
rect 17221 10047 17279 10053
rect 17221 10044 17233 10047
rect 17184 10016 17233 10044
rect 17184 10004 17190 10016
rect 17221 10013 17233 10016
rect 17267 10013 17279 10047
rect 17221 10007 17279 10013
rect 15580 9976 15608 10004
rect 16669 9979 16727 9985
rect 16669 9976 16681 9979
rect 14844 9948 16681 9976
rect 16669 9945 16681 9948
rect 16715 9945 16727 9979
rect 16669 9939 16727 9945
rect 2556 9880 6592 9908
rect 2556 9868 2562 9880
rect 10042 9868 10048 9920
rect 10100 9908 10106 9920
rect 10962 9908 10968 9920
rect 10100 9880 10968 9908
rect 10100 9868 10106 9880
rect 10962 9868 10968 9880
rect 11020 9868 11026 9920
rect 12437 9911 12495 9917
rect 12437 9877 12449 9911
rect 12483 9908 12495 9911
rect 12526 9908 12532 9920
rect 12483 9880 12532 9908
rect 12483 9877 12495 9880
rect 12437 9871 12495 9877
rect 12526 9868 12532 9880
rect 12584 9868 12590 9920
rect 12710 9868 12716 9920
rect 12768 9868 12774 9920
rect 12894 9868 12900 9920
rect 12952 9868 12958 9920
rect 14550 9868 14556 9920
rect 14608 9908 14614 9920
rect 14737 9911 14795 9917
rect 14737 9908 14749 9911
rect 14608 9880 14749 9908
rect 14608 9868 14614 9880
rect 14737 9877 14749 9880
rect 14783 9877 14795 9911
rect 14737 9871 14795 9877
rect 15197 9911 15255 9917
rect 15197 9877 15209 9911
rect 15243 9908 15255 9911
rect 15562 9908 15568 9920
rect 15243 9880 15568 9908
rect 15243 9877 15255 9880
rect 15197 9871 15255 9877
rect 15562 9868 15568 9880
rect 15620 9868 15626 9920
rect 16574 9868 16580 9920
rect 16632 9868 16638 9920
rect 16853 9911 16911 9917
rect 16853 9877 16865 9911
rect 16899 9908 16911 9911
rect 17129 9911 17187 9917
rect 17129 9908 17141 9911
rect 16899 9880 17141 9908
rect 16899 9877 16911 9880
rect 16853 9871 16911 9877
rect 17129 9877 17141 9880
rect 17175 9877 17187 9911
rect 17129 9871 17187 9877
rect 1104 9818 17848 9840
rect 1104 9766 2658 9818
rect 2710 9766 2722 9818
rect 2774 9766 2786 9818
rect 2838 9766 2850 9818
rect 2902 9766 2914 9818
rect 2966 9766 2978 9818
rect 3030 9766 8658 9818
rect 8710 9766 8722 9818
rect 8774 9766 8786 9818
rect 8838 9766 8850 9818
rect 8902 9766 8914 9818
rect 8966 9766 8978 9818
rect 9030 9766 14658 9818
rect 14710 9766 14722 9818
rect 14774 9766 14786 9818
rect 14838 9766 14850 9818
rect 14902 9766 14914 9818
rect 14966 9766 14978 9818
rect 15030 9766 17848 9818
rect 1104 9744 17848 9766
rect 3237 9707 3295 9713
rect 3237 9673 3249 9707
rect 3283 9704 3295 9707
rect 3878 9704 3884 9716
rect 3283 9676 3884 9704
rect 3283 9673 3295 9676
rect 3237 9667 3295 9673
rect 3878 9664 3884 9676
rect 3936 9664 3942 9716
rect 4525 9707 4583 9713
rect 4525 9704 4537 9707
rect 4264 9676 4537 9704
rect 2406 9596 2412 9648
rect 2464 9596 2470 9648
rect 3605 9639 3663 9645
rect 3605 9605 3617 9639
rect 3651 9636 3663 9639
rect 4264 9636 4292 9676
rect 4525 9673 4537 9676
rect 4571 9673 4583 9707
rect 4525 9667 4583 9673
rect 5077 9707 5135 9713
rect 5077 9673 5089 9707
rect 5123 9673 5135 9707
rect 5077 9667 5135 9673
rect 10137 9707 10195 9713
rect 10137 9673 10149 9707
rect 10183 9673 10195 9707
rect 12618 9704 12624 9716
rect 10137 9667 10195 9673
rect 11992 9676 12624 9704
rect 5092 9636 5120 9667
rect 3651 9608 4292 9636
rect 3651 9605 3663 9608
rect 3605 9599 3663 9605
rect 1394 9528 1400 9580
rect 1452 9568 1458 9580
rect 1581 9571 1639 9577
rect 1581 9568 1593 9571
rect 1452 9540 1593 9568
rect 1452 9528 1458 9540
rect 1581 9537 1593 9540
rect 1627 9537 1639 9571
rect 2498 9568 2504 9580
rect 1581 9531 1639 9537
rect 2424 9540 2504 9568
rect 2424 9512 2452 9540
rect 2498 9528 2504 9540
rect 2556 9528 2562 9580
rect 3418 9528 3424 9580
rect 3476 9528 3482 9580
rect 3510 9528 3516 9580
rect 3568 9528 3574 9580
rect 3789 9571 3847 9577
rect 3789 9537 3801 9571
rect 3835 9568 3847 9571
rect 3970 9568 3976 9580
rect 3835 9540 3976 9568
rect 3835 9537 3847 9540
rect 3789 9531 3847 9537
rect 3970 9528 3976 9540
rect 4028 9528 4034 9580
rect 4062 9528 4068 9580
rect 4120 9568 4126 9580
rect 4264 9568 4292 9608
rect 4356 9608 5120 9636
rect 5245 9639 5303 9645
rect 4356 9577 4384 9608
rect 5245 9605 5257 9639
rect 5291 9636 5303 9639
rect 5445 9639 5503 9645
rect 5291 9605 5304 9636
rect 5245 9599 5304 9605
rect 5445 9605 5457 9639
rect 5491 9636 5503 9639
rect 5718 9636 5724 9648
rect 5491 9608 5724 9636
rect 5491 9605 5503 9608
rect 5445 9599 5503 9605
rect 4120 9540 4292 9568
rect 4341 9571 4399 9577
rect 4120 9528 4126 9540
rect 4341 9537 4353 9571
rect 4387 9537 4399 9571
rect 4341 9531 4399 9537
rect 4706 9528 4712 9580
rect 4764 9528 4770 9580
rect 4890 9528 4896 9580
rect 4948 9528 4954 9580
rect 4985 9571 5043 9577
rect 4985 9537 4997 9571
rect 5031 9568 5043 9571
rect 5074 9568 5080 9580
rect 5031 9540 5080 9568
rect 5031 9537 5043 9540
rect 4985 9531 5043 9537
rect 5074 9528 5080 9540
rect 5132 9528 5138 9580
rect 2406 9460 2412 9512
rect 2464 9460 2470 9512
rect 3694 9460 3700 9512
rect 3752 9500 3758 9512
rect 3881 9503 3939 9509
rect 3881 9500 3893 9503
rect 3752 9472 3893 9500
rect 3752 9460 3758 9472
rect 3881 9469 3893 9472
rect 3927 9469 3939 9503
rect 3881 9463 3939 9469
rect 4154 9460 4160 9512
rect 4212 9460 4218 9512
rect 4249 9503 4307 9509
rect 4249 9469 4261 9503
rect 4295 9500 4307 9503
rect 4430 9500 4436 9512
rect 4295 9472 4436 9500
rect 4295 9469 4307 9472
rect 4249 9463 4307 9469
rect 4430 9460 4436 9472
rect 4488 9460 4494 9512
rect 4724 9500 4752 9528
rect 5276 9500 5304 9599
rect 5718 9596 5724 9608
rect 5776 9596 5782 9648
rect 8113 9639 8171 9645
rect 8113 9605 8125 9639
rect 8159 9636 8171 9639
rect 9674 9636 9680 9648
rect 8159 9608 9680 9636
rect 8159 9605 8171 9608
rect 8113 9599 8171 9605
rect 9674 9596 9680 9608
rect 9732 9596 9738 9648
rect 10152 9636 10180 9667
rect 10152 9608 10548 9636
rect 5813 9571 5871 9577
rect 5813 9537 5825 9571
rect 5859 9568 5871 9571
rect 6365 9571 6423 9577
rect 6365 9568 6377 9571
rect 5859 9540 6377 9568
rect 5859 9537 5871 9540
rect 5813 9531 5871 9537
rect 6365 9537 6377 9540
rect 6411 9537 6423 9571
rect 6365 9531 6423 9537
rect 8757 9571 8815 9577
rect 8757 9537 8769 9571
rect 8803 9568 8815 9571
rect 9217 9571 9275 9577
rect 9217 9568 9229 9571
rect 8803 9540 9229 9568
rect 8803 9537 8815 9540
rect 8757 9531 8815 9537
rect 9217 9537 9229 9540
rect 9263 9568 9275 9571
rect 9263 9540 9720 9568
rect 9263 9537 9275 9540
rect 9217 9531 9275 9537
rect 4724 9472 5304 9500
rect 1302 9392 1308 9444
rect 1360 9432 1366 9444
rect 1397 9435 1455 9441
rect 1397 9432 1409 9435
rect 1360 9404 1409 9432
rect 1360 9392 1366 9404
rect 1397 9401 1409 9404
rect 1443 9401 1455 9435
rect 1397 9395 1455 9401
rect 3142 9392 3148 9444
rect 3200 9432 3206 9444
rect 5828 9432 5856 9531
rect 8386 9460 8392 9512
rect 8444 9500 8450 9512
rect 8665 9503 8723 9509
rect 8665 9500 8677 9503
rect 8444 9472 8677 9500
rect 8444 9460 8450 9472
rect 8665 9469 8677 9472
rect 8711 9469 8723 9503
rect 8665 9463 8723 9469
rect 9493 9503 9551 9509
rect 9493 9469 9505 9503
rect 9539 9469 9551 9503
rect 9493 9463 9551 9469
rect 3200 9404 5856 9432
rect 3200 9392 3206 9404
rect 9508 9376 9536 9463
rect 9692 9432 9720 9540
rect 9766 9528 9772 9580
rect 9824 9528 9830 9580
rect 9861 9503 9919 9509
rect 9861 9469 9873 9503
rect 9907 9500 9919 9503
rect 10042 9500 10048 9512
rect 9907 9472 10048 9500
rect 9907 9469 9919 9472
rect 9861 9463 9919 9469
rect 10042 9460 10048 9472
rect 10100 9460 10106 9512
rect 10520 9509 10548 9608
rect 10597 9571 10655 9577
rect 10597 9537 10609 9571
rect 10643 9568 10655 9571
rect 10686 9568 10692 9580
rect 10643 9540 10692 9568
rect 10643 9537 10655 9540
rect 10597 9531 10655 9537
rect 10686 9528 10692 9540
rect 10744 9528 10750 9580
rect 11330 9528 11336 9580
rect 11388 9568 11394 9580
rect 11701 9571 11759 9577
rect 11701 9568 11713 9571
rect 11388 9540 11713 9568
rect 11388 9528 11394 9540
rect 11701 9537 11713 9540
rect 11747 9537 11759 9571
rect 11701 9531 11759 9537
rect 11793 9571 11851 9577
rect 11793 9537 11805 9571
rect 11839 9568 11851 9571
rect 11992 9568 12020 9676
rect 12618 9664 12624 9676
rect 12676 9704 12682 9716
rect 13078 9704 13084 9716
rect 12676 9676 13084 9704
rect 12676 9664 12682 9676
rect 13078 9664 13084 9676
rect 13136 9664 13142 9716
rect 15470 9704 15476 9716
rect 14476 9676 15476 9704
rect 13725 9639 13783 9645
rect 13725 9636 13737 9639
rect 11839 9540 12020 9568
rect 12176 9608 13737 9636
rect 11839 9537 11851 9540
rect 11793 9531 11851 9537
rect 10505 9503 10563 9509
rect 10505 9469 10517 9503
rect 10551 9469 10563 9503
rect 10505 9463 10563 9469
rect 11974 9460 11980 9512
rect 12032 9460 12038 9512
rect 12176 9432 12204 9608
rect 13725 9605 13737 9608
rect 13771 9605 13783 9639
rect 13725 9599 13783 9605
rect 14182 9596 14188 9648
rect 14240 9596 14246 9648
rect 12253 9571 12311 9577
rect 12253 9537 12265 9571
rect 12299 9537 12311 9571
rect 12253 9531 12311 9537
rect 12345 9571 12403 9577
rect 12345 9537 12357 9571
rect 12391 9537 12403 9571
rect 12345 9531 12403 9537
rect 9692 9404 12204 9432
rect 3418 9324 3424 9376
rect 3476 9364 3482 9376
rect 4154 9364 4160 9376
rect 3476 9336 4160 9364
rect 3476 9324 3482 9336
rect 4154 9324 4160 9336
rect 4212 9324 4218 9376
rect 5258 9324 5264 9376
rect 5316 9324 5322 9376
rect 7282 9324 7288 9376
rect 7340 9364 7346 9376
rect 8481 9367 8539 9373
rect 8481 9364 8493 9367
rect 7340 9336 8493 9364
rect 7340 9324 7346 9336
rect 8481 9333 8493 9336
rect 8527 9333 8539 9367
rect 8481 9327 8539 9333
rect 8662 9324 8668 9376
rect 8720 9364 8726 9376
rect 9033 9367 9091 9373
rect 9033 9364 9045 9367
rect 8720 9336 9045 9364
rect 8720 9324 8726 9336
rect 9033 9333 9045 9336
rect 9079 9333 9091 9367
rect 9033 9327 9091 9333
rect 9214 9324 9220 9376
rect 9272 9364 9278 9376
rect 9401 9367 9459 9373
rect 9401 9364 9413 9367
rect 9272 9336 9413 9364
rect 9272 9324 9278 9336
rect 9401 9333 9413 9336
rect 9447 9333 9459 9367
rect 9401 9327 9459 9333
rect 9490 9324 9496 9376
rect 9548 9364 9554 9376
rect 10321 9367 10379 9373
rect 10321 9364 10333 9367
rect 9548 9336 10333 9364
rect 9548 9324 9554 9336
rect 10321 9333 10333 9336
rect 10367 9333 10379 9367
rect 10321 9327 10379 9333
rect 11882 9324 11888 9376
rect 11940 9324 11946 9376
rect 12066 9324 12072 9376
rect 12124 9324 12130 9376
rect 12268 9364 12296 9531
rect 12360 9500 12388 9531
rect 12526 9528 12532 9580
rect 12584 9528 12590 9580
rect 12618 9528 12624 9580
rect 12676 9528 12682 9580
rect 12894 9528 12900 9580
rect 12952 9528 12958 9580
rect 13078 9528 13084 9580
rect 13136 9528 13142 9580
rect 13446 9528 13452 9580
rect 13504 9528 13510 9580
rect 13814 9528 13820 9580
rect 13872 9568 13878 9580
rect 13909 9571 13967 9577
rect 13909 9568 13921 9571
rect 13872 9540 13921 9568
rect 13872 9528 13878 9540
rect 13909 9537 13921 9540
rect 13955 9537 13967 9571
rect 13909 9531 13967 9537
rect 14001 9571 14059 9577
rect 14001 9537 14013 9571
rect 14047 9537 14059 9571
rect 14200 9568 14228 9596
rect 14277 9571 14335 9577
rect 14277 9568 14289 9571
rect 14200 9540 14289 9568
rect 14001 9531 14059 9537
rect 14277 9537 14289 9540
rect 14323 9537 14335 9571
rect 14476 9574 14504 9676
rect 15470 9664 15476 9676
rect 15528 9664 15534 9716
rect 15194 9636 15200 9648
rect 15028 9608 15200 9636
rect 14553 9574 14611 9577
rect 14476 9571 14611 9574
rect 14476 9546 14565 9571
rect 14277 9531 14335 9537
rect 14553 9537 14565 9546
rect 14599 9537 14611 9571
rect 14553 9531 14611 9537
rect 14737 9571 14795 9577
rect 14737 9537 14749 9571
rect 14783 9568 14795 9571
rect 14918 9568 14924 9580
rect 14783 9540 14924 9568
rect 14783 9537 14795 9540
rect 14737 9531 14795 9537
rect 12986 9500 12992 9512
rect 12360 9472 12992 9500
rect 12986 9460 12992 9472
rect 13044 9460 13050 9512
rect 13170 9460 13176 9512
rect 13228 9460 13234 9512
rect 13265 9503 13323 9509
rect 13265 9469 13277 9503
rect 13311 9469 13323 9503
rect 13265 9463 13323 9469
rect 13633 9503 13691 9509
rect 13633 9469 13645 9503
rect 13679 9500 13691 9503
rect 13725 9503 13783 9509
rect 13725 9500 13737 9503
rect 13679 9472 13737 9500
rect 13679 9469 13691 9472
rect 13633 9463 13691 9469
rect 13725 9469 13737 9472
rect 13771 9469 13783 9503
rect 14016 9500 14044 9531
rect 14918 9528 14924 9540
rect 14976 9528 14982 9580
rect 15028 9577 15056 9608
rect 15194 9596 15200 9608
rect 15252 9596 15258 9648
rect 16114 9636 16120 9648
rect 15488 9608 15700 9636
rect 15378 9583 15384 9586
rect 15013 9571 15071 9577
rect 15377 9574 15384 9583
rect 15013 9537 15025 9571
rect 15059 9537 15071 9571
rect 15304 9568 15384 9574
rect 15013 9531 15071 9537
rect 15120 9546 15384 9568
rect 15120 9540 15332 9546
rect 15120 9512 15148 9540
rect 15377 9537 15384 9546
rect 15378 9534 15384 9537
rect 15436 9534 15442 9586
rect 15488 9580 15516 9608
rect 15672 9580 15700 9608
rect 15856 9608 16120 9636
rect 15470 9528 15476 9580
rect 15528 9528 15534 9580
rect 15562 9528 15568 9580
rect 15620 9528 15626 9580
rect 15654 9528 15660 9580
rect 15712 9528 15718 9580
rect 15746 9528 15752 9580
rect 15804 9528 15810 9580
rect 15856 9577 15884 9608
rect 16114 9596 16120 9608
rect 16172 9636 16178 9648
rect 16172 9608 17080 9636
rect 16172 9596 16178 9608
rect 15841 9571 15899 9577
rect 15841 9537 15853 9571
rect 15887 9537 15899 9571
rect 15841 9531 15899 9537
rect 16574 9528 16580 9580
rect 16632 9568 16638 9580
rect 16669 9571 16727 9577
rect 16669 9568 16681 9571
rect 16632 9540 16681 9568
rect 16632 9528 16638 9540
rect 16669 9537 16681 9540
rect 16715 9537 16727 9571
rect 16669 9531 16727 9537
rect 16850 9528 16856 9580
rect 16908 9528 16914 9580
rect 17052 9577 17080 9608
rect 17037 9571 17095 9577
rect 17037 9537 17049 9571
rect 17083 9537 17095 9571
rect 17037 9531 17095 9537
rect 17218 9528 17224 9580
rect 17276 9528 17282 9580
rect 14016 9472 14228 9500
rect 13725 9463 13783 9469
rect 12802 9392 12808 9444
rect 12860 9432 12866 9444
rect 13280 9432 13308 9463
rect 12860 9404 13308 9432
rect 12860 9392 12866 9404
rect 13354 9392 13360 9444
rect 13412 9432 13418 9444
rect 14093 9435 14151 9441
rect 14093 9432 14105 9435
rect 13412 9404 14105 9432
rect 13412 9392 13418 9404
rect 14093 9401 14105 9404
rect 14139 9401 14151 9435
rect 14093 9395 14151 9401
rect 12434 9364 12440 9376
rect 12268 9336 12440 9364
rect 12434 9324 12440 9336
rect 12492 9324 12498 9376
rect 13446 9324 13452 9376
rect 13504 9364 13510 9376
rect 13998 9364 14004 9376
rect 13504 9336 14004 9364
rect 13504 9324 13510 9336
rect 13998 9324 14004 9336
rect 14056 9324 14062 9376
rect 14200 9364 14228 9472
rect 14458 9460 14464 9512
rect 14516 9460 14522 9512
rect 15102 9460 15108 9512
rect 15160 9460 15166 9512
rect 15197 9503 15255 9509
rect 15197 9469 15209 9503
rect 15243 9469 15255 9503
rect 15197 9463 15255 9469
rect 14369 9435 14427 9441
rect 14369 9401 14381 9435
rect 14415 9432 14427 9435
rect 14918 9432 14924 9444
rect 14415 9404 14924 9432
rect 14415 9401 14427 9404
rect 14369 9395 14427 9401
rect 14918 9392 14924 9404
rect 14976 9392 14982 9444
rect 14550 9364 14556 9376
rect 14200 9336 14556 9364
rect 14550 9324 14556 9336
rect 14608 9324 14614 9376
rect 14829 9367 14887 9373
rect 14829 9333 14841 9367
rect 14875 9364 14887 9367
rect 15010 9364 15016 9376
rect 14875 9336 15016 9364
rect 14875 9333 14887 9336
rect 14829 9327 14887 9333
rect 15010 9324 15016 9336
rect 15068 9324 15074 9376
rect 15212 9364 15240 9463
rect 15286 9460 15292 9512
rect 15344 9460 15350 9512
rect 16945 9503 17003 9509
rect 16945 9469 16957 9503
rect 16991 9500 17003 9503
rect 17126 9500 17132 9512
rect 16991 9472 17132 9500
rect 16991 9469 17003 9472
rect 16945 9463 17003 9469
rect 17126 9460 17132 9472
rect 17184 9460 17190 9512
rect 16114 9364 16120 9376
rect 15212 9336 16120 9364
rect 16114 9324 16120 9336
rect 16172 9324 16178 9376
rect 17034 9324 17040 9376
rect 17092 9364 17098 9376
rect 17405 9367 17463 9373
rect 17405 9364 17417 9367
rect 17092 9336 17417 9364
rect 17092 9324 17098 9336
rect 17405 9333 17417 9336
rect 17451 9333 17463 9367
rect 17405 9327 17463 9333
rect 1104 9274 17848 9296
rect 1104 9222 1918 9274
rect 1970 9222 1982 9274
rect 2034 9222 2046 9274
rect 2098 9222 2110 9274
rect 2162 9222 2174 9274
rect 2226 9222 2238 9274
rect 2290 9222 7918 9274
rect 7970 9222 7982 9274
rect 8034 9222 8046 9274
rect 8098 9222 8110 9274
rect 8162 9222 8174 9274
rect 8226 9222 8238 9274
rect 8290 9222 13918 9274
rect 13970 9222 13982 9274
rect 14034 9222 14046 9274
rect 14098 9222 14110 9274
rect 14162 9222 14174 9274
rect 14226 9222 14238 9274
rect 14290 9222 17848 9274
rect 1104 9200 17848 9222
rect 1394 9120 1400 9172
rect 1452 9120 1458 9172
rect 3510 9120 3516 9172
rect 3568 9160 3574 9172
rect 4154 9160 4160 9172
rect 3568 9132 4160 9160
rect 3568 9120 3574 9132
rect 3804 9101 3832 9132
rect 4154 9120 4160 9132
rect 4212 9120 4218 9172
rect 4246 9120 4252 9172
rect 4304 9160 4310 9172
rect 4341 9163 4399 9169
rect 4341 9160 4353 9163
rect 4304 9132 4353 9160
rect 4304 9120 4310 9132
rect 4341 9129 4353 9132
rect 4387 9129 4399 9163
rect 4341 9123 4399 9129
rect 6914 9120 6920 9172
rect 6972 9160 6978 9172
rect 7101 9163 7159 9169
rect 7101 9160 7113 9163
rect 6972 9132 7113 9160
rect 6972 9120 6978 9132
rect 7101 9129 7113 9132
rect 7147 9129 7159 9163
rect 7101 9123 7159 9129
rect 8297 9163 8355 9169
rect 8297 9129 8309 9163
rect 8343 9160 8355 9163
rect 8386 9160 8392 9172
rect 8343 9132 8392 9160
rect 8343 9129 8355 9132
rect 8297 9123 8355 9129
rect 8386 9120 8392 9132
rect 8444 9120 8450 9172
rect 8478 9120 8484 9172
rect 8536 9160 8542 9172
rect 8665 9163 8723 9169
rect 8665 9160 8677 9163
rect 8536 9132 8677 9160
rect 8536 9120 8542 9132
rect 8665 9129 8677 9132
rect 8711 9129 8723 9163
rect 12066 9160 12072 9172
rect 8665 9123 8723 9129
rect 8772 9132 12072 9160
rect 3789 9095 3847 9101
rect 3789 9061 3801 9095
rect 3835 9061 3847 9095
rect 4617 9095 4675 9101
rect 4617 9092 4629 9095
rect 3789 9055 3847 9061
rect 4172 9064 4629 9092
rect 3142 8984 3148 9036
rect 3200 8984 3206 9036
rect 3970 8916 3976 8968
rect 4028 8956 4034 8968
rect 4172 8965 4200 9064
rect 4617 9061 4629 9064
rect 4663 9061 4675 9095
rect 8772 9092 8800 9132
rect 12066 9120 12072 9132
rect 12124 9120 12130 9172
rect 12618 9120 12624 9172
rect 12676 9120 12682 9172
rect 14369 9163 14427 9169
rect 14369 9129 14381 9163
rect 14415 9160 14427 9163
rect 14550 9160 14556 9172
rect 14415 9132 14556 9160
rect 14415 9129 14427 9132
rect 14369 9123 14427 9129
rect 14550 9120 14556 9132
rect 14608 9120 14614 9172
rect 14918 9120 14924 9172
rect 14976 9160 14982 9172
rect 15105 9163 15163 9169
rect 15105 9160 15117 9163
rect 14976 9132 15117 9160
rect 14976 9120 14982 9132
rect 15105 9129 15117 9132
rect 15151 9129 15163 9163
rect 15105 9123 15163 9129
rect 4617 9055 4675 9061
rect 6656 9064 8800 9092
rect 4706 9024 4712 9036
rect 4540 8996 4712 9024
rect 4540 8965 4568 8996
rect 4706 8984 4712 8996
rect 4764 9024 4770 9036
rect 6457 9027 6515 9033
rect 6457 9024 6469 9027
rect 4764 8996 6469 9024
rect 4764 8984 4770 8996
rect 6457 8993 6469 8996
rect 6503 8993 6515 9027
rect 6457 8987 6515 8993
rect 4157 8959 4215 8965
rect 4157 8956 4169 8959
rect 4028 8928 4169 8956
rect 4028 8916 4034 8928
rect 4157 8925 4169 8928
rect 4203 8925 4215 8959
rect 4157 8919 4215 8925
rect 4525 8959 4583 8965
rect 4525 8925 4537 8959
rect 4571 8925 4583 8959
rect 4525 8919 4583 8925
rect 4801 8959 4859 8965
rect 4801 8925 4813 8959
rect 4847 8956 4859 8959
rect 4890 8956 4896 8968
rect 4847 8928 4896 8956
rect 4847 8925 4859 8928
rect 4801 8919 4859 8925
rect 4890 8916 4896 8928
rect 4948 8956 4954 8968
rect 4948 8928 5396 8956
rect 4948 8916 4954 8928
rect 2222 8848 2228 8900
rect 2280 8848 2286 8900
rect 2869 8891 2927 8897
rect 2869 8857 2881 8891
rect 2915 8857 2927 8891
rect 2869 8851 2927 8857
rect 2884 8820 2912 8851
rect 4062 8848 4068 8900
rect 4120 8848 4126 8900
rect 4709 8891 4767 8897
rect 4709 8857 4721 8891
rect 4755 8888 4767 8891
rect 5258 8888 5264 8900
rect 4755 8860 5264 8888
rect 4755 8857 4767 8860
rect 4709 8851 4767 8857
rect 5258 8848 5264 8860
rect 5316 8848 5322 8900
rect 5368 8888 5396 8928
rect 5534 8916 5540 8968
rect 5592 8916 5598 8968
rect 5626 8916 5632 8968
rect 5684 8956 5690 8968
rect 5997 8959 6055 8965
rect 5997 8956 6009 8959
rect 5684 8928 6009 8956
rect 5684 8916 5690 8928
rect 5997 8925 6009 8928
rect 6043 8956 6055 8959
rect 6656 8956 6684 9064
rect 9674 9052 9680 9104
rect 9732 9092 9738 9104
rect 13354 9092 13360 9104
rect 9732 9064 13360 9092
rect 9732 9052 9738 9064
rect 13354 9052 13360 9064
rect 13412 9052 13418 9104
rect 15194 9092 15200 9104
rect 14384 9064 15200 9092
rect 6733 9027 6791 9033
rect 6733 8993 6745 9027
rect 6779 8993 6791 9027
rect 8021 9027 8079 9033
rect 6733 8987 6791 8993
rect 6840 8996 7328 9024
rect 6043 8928 6684 8956
rect 6043 8925 6055 8928
rect 5997 8919 6055 8925
rect 5718 8888 5724 8900
rect 5368 8860 5724 8888
rect 5718 8848 5724 8860
rect 5776 8848 5782 8900
rect 6748 8888 6776 8987
rect 6840 8965 6868 8996
rect 7300 8968 7328 8996
rect 8021 8993 8033 9027
rect 8067 9024 8079 9027
rect 9214 9024 9220 9036
rect 8067 8996 9220 9024
rect 8067 8993 8079 8996
rect 8021 8987 8079 8993
rect 6825 8959 6883 8965
rect 6825 8925 6837 8959
rect 6871 8925 6883 8959
rect 6825 8919 6883 8925
rect 7101 8959 7159 8965
rect 7101 8925 7113 8959
rect 7147 8925 7159 8959
rect 7101 8919 7159 8925
rect 7116 8888 7144 8919
rect 7282 8916 7288 8968
rect 7340 8916 7346 8968
rect 8404 8965 8432 8996
rect 9214 8984 9220 8996
rect 9272 8984 9278 9036
rect 11974 8984 11980 9036
rect 12032 9024 12038 9036
rect 12802 9024 12808 9036
rect 12032 8996 12808 9024
rect 12032 8984 12038 8996
rect 7929 8959 7987 8965
rect 7929 8925 7941 8959
rect 7975 8925 7987 8959
rect 7929 8919 7987 8925
rect 8389 8959 8447 8965
rect 8389 8925 8401 8959
rect 8435 8925 8447 8959
rect 8389 8919 8447 8925
rect 7374 8888 7380 8900
rect 6748 8860 7380 8888
rect 7374 8848 7380 8860
rect 7432 8848 7438 8900
rect 7944 8888 7972 8919
rect 8662 8916 8668 8968
rect 8720 8916 8726 8968
rect 12360 8965 12388 8996
rect 12802 8984 12808 8996
rect 12860 8984 12866 9036
rect 12345 8959 12403 8965
rect 12345 8925 12357 8959
rect 12391 8925 12403 8959
rect 12345 8919 12403 8925
rect 12621 8959 12679 8965
rect 12621 8925 12633 8959
rect 12667 8956 12679 8959
rect 12710 8956 12716 8968
rect 12667 8928 12716 8956
rect 12667 8925 12679 8928
rect 12621 8919 12679 8925
rect 12710 8916 12716 8928
rect 12768 8916 12774 8968
rect 13170 8916 13176 8968
rect 13228 8956 13234 8968
rect 14277 8959 14335 8965
rect 14277 8956 14289 8959
rect 13228 8928 14289 8956
rect 13228 8916 13234 8928
rect 14277 8925 14289 8928
rect 14323 8956 14335 8959
rect 14384 8956 14412 9064
rect 15194 9052 15200 9064
rect 15252 9052 15258 9104
rect 15286 9052 15292 9104
rect 15344 9092 15350 9104
rect 17218 9092 17224 9104
rect 15344 9064 17224 9092
rect 15344 9052 15350 9064
rect 14458 8984 14464 9036
rect 14516 9024 14522 9036
rect 16684 9033 16712 9064
rect 17218 9052 17224 9064
rect 17276 9052 17282 9104
rect 16577 9027 16635 9033
rect 16577 9024 16589 9027
rect 14516 8996 16589 9024
rect 14516 8984 14522 8996
rect 14752 8965 14780 8996
rect 16577 8993 16589 8996
rect 16623 8993 16635 9027
rect 16577 8987 16635 8993
rect 16669 9027 16727 9033
rect 16669 8993 16681 9027
rect 16715 8993 16727 9027
rect 16669 8987 16727 8993
rect 17034 8984 17040 9036
rect 17092 8984 17098 9036
rect 14323 8928 14412 8956
rect 14737 8959 14795 8965
rect 14323 8925 14335 8928
rect 14277 8919 14335 8925
rect 14737 8925 14749 8959
rect 14783 8925 14795 8959
rect 14737 8919 14795 8925
rect 15010 8916 15016 8968
rect 15068 8916 15074 8968
rect 15102 8916 15108 8968
rect 15160 8916 15166 8968
rect 15194 8916 15200 8968
rect 15252 8956 15258 8968
rect 15289 8959 15347 8965
rect 15289 8956 15301 8959
rect 15252 8928 15301 8956
rect 15252 8916 15258 8928
rect 15289 8925 15301 8928
rect 15335 8956 15347 8959
rect 15838 8956 15844 8968
rect 15335 8928 15844 8956
rect 15335 8925 15347 8928
rect 15289 8919 15347 8925
rect 15838 8916 15844 8928
rect 15896 8916 15902 8968
rect 16850 8956 16856 8968
rect 15948 8928 16856 8956
rect 8481 8891 8539 8897
rect 8481 8888 8493 8891
rect 7944 8860 8493 8888
rect 8481 8857 8493 8860
rect 8527 8888 8539 8891
rect 9490 8888 9496 8900
rect 8527 8860 9496 8888
rect 8527 8857 8539 8860
rect 8481 8851 8539 8857
rect 9490 8848 9496 8860
rect 9548 8848 9554 8900
rect 14550 8848 14556 8900
rect 14608 8888 14614 8900
rect 14829 8891 14887 8897
rect 14829 8888 14841 8891
rect 14608 8860 14841 8888
rect 14608 8848 14614 8860
rect 14829 8857 14841 8860
rect 14875 8857 14887 8891
rect 15120 8888 15148 8916
rect 15948 8888 15976 8928
rect 16850 8916 16856 8928
rect 16908 8916 16914 8968
rect 17126 8916 17132 8968
rect 17184 8916 17190 8968
rect 15120 8860 15976 8888
rect 14829 8851 14887 8857
rect 16758 8848 16764 8900
rect 16816 8888 16822 8900
rect 17221 8891 17279 8897
rect 17221 8888 17233 8891
rect 16816 8860 17233 8888
rect 16816 8848 16822 8860
rect 17221 8857 17233 8860
rect 17267 8857 17279 8891
rect 17221 8851 17279 8857
rect 3050 8820 3056 8832
rect 2884 8792 3056 8820
rect 3050 8780 3056 8792
rect 3108 8780 3114 8832
rect 3970 8780 3976 8832
rect 4028 8820 4034 8832
rect 5169 8823 5227 8829
rect 5169 8820 5181 8823
rect 4028 8792 5181 8820
rect 4028 8780 4034 8792
rect 5169 8789 5181 8792
rect 5215 8789 5227 8823
rect 5169 8783 5227 8789
rect 12437 8823 12495 8829
rect 12437 8789 12449 8823
rect 12483 8820 12495 8823
rect 12710 8820 12716 8832
rect 12483 8792 12716 8820
rect 12483 8789 12495 8792
rect 12437 8783 12495 8789
rect 12710 8780 12716 8792
rect 12768 8820 12774 8832
rect 13262 8820 13268 8832
rect 12768 8792 13268 8820
rect 12768 8780 12774 8792
rect 13262 8780 13268 8792
rect 13320 8780 13326 8832
rect 14914 8823 14972 8829
rect 14914 8789 14926 8823
rect 14960 8820 14972 8823
rect 15102 8820 15108 8832
rect 14960 8792 15108 8820
rect 14960 8789 14972 8792
rect 14914 8783 14972 8789
rect 15102 8780 15108 8792
rect 15160 8780 15166 8832
rect 16390 8780 16396 8832
rect 16448 8780 16454 8832
rect 1104 8730 17848 8752
rect 1104 8678 2658 8730
rect 2710 8678 2722 8730
rect 2774 8678 2786 8730
rect 2838 8678 2850 8730
rect 2902 8678 2914 8730
rect 2966 8678 2978 8730
rect 3030 8678 8658 8730
rect 8710 8678 8722 8730
rect 8774 8678 8786 8730
rect 8838 8678 8850 8730
rect 8902 8678 8914 8730
rect 8966 8678 8978 8730
rect 9030 8678 14658 8730
rect 14710 8678 14722 8730
rect 14774 8678 14786 8730
rect 14838 8678 14850 8730
rect 14902 8678 14914 8730
rect 14966 8678 14978 8730
rect 15030 8678 17848 8730
rect 1104 8656 17848 8678
rect 1302 8576 1308 8628
rect 1360 8616 1366 8628
rect 1397 8619 1455 8625
rect 1397 8616 1409 8619
rect 1360 8588 1409 8616
rect 1360 8576 1366 8588
rect 1397 8585 1409 8588
rect 1443 8585 1455 8619
rect 1397 8579 1455 8585
rect 2222 8576 2228 8628
rect 2280 8576 2286 8628
rect 5258 8576 5264 8628
rect 5316 8616 5322 8628
rect 5445 8619 5503 8625
rect 5445 8616 5457 8619
rect 5316 8588 5457 8616
rect 5316 8576 5322 8588
rect 5445 8585 5457 8588
rect 5491 8585 5503 8619
rect 5445 8579 5503 8585
rect 5718 8576 5724 8628
rect 5776 8576 5782 8628
rect 9214 8576 9220 8628
rect 9272 8576 9278 8628
rect 11514 8576 11520 8628
rect 11572 8616 11578 8628
rect 12069 8619 12127 8625
rect 12069 8616 12081 8619
rect 11572 8588 12081 8616
rect 11572 8576 11578 8588
rect 12069 8585 12081 8588
rect 12115 8585 12127 8619
rect 17126 8616 17132 8628
rect 12069 8579 12127 8585
rect 12406 8588 17132 8616
rect 11882 8548 11888 8560
rect 5368 8520 5948 8548
rect 5368 8492 5396 8520
rect 1578 8440 1584 8492
rect 1636 8440 1642 8492
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8480 2191 8483
rect 2406 8480 2412 8492
rect 2179 8452 2412 8480
rect 2179 8449 2191 8452
rect 2133 8443 2191 8449
rect 2406 8440 2412 8452
rect 2464 8440 2470 8492
rect 3237 8483 3295 8489
rect 3237 8449 3249 8483
rect 3283 8480 3295 8483
rect 4154 8480 4160 8492
rect 3283 8452 4160 8480
rect 3283 8449 3295 8452
rect 3237 8443 3295 8449
rect 4154 8440 4160 8452
rect 4212 8440 4218 8492
rect 5166 8440 5172 8492
rect 5224 8489 5230 8492
rect 5224 8483 5246 8489
rect 5234 8449 5246 8483
rect 5224 8443 5246 8449
rect 5224 8440 5230 8443
rect 5350 8440 5356 8492
rect 5408 8440 5414 8492
rect 5626 8440 5632 8492
rect 5684 8440 5690 8492
rect 5920 8489 5948 8520
rect 7760 8520 11888 8548
rect 5721 8483 5779 8489
rect 5721 8449 5733 8483
rect 5767 8449 5779 8483
rect 5721 8443 5779 8449
rect 5905 8483 5963 8489
rect 5905 8449 5917 8483
rect 5951 8480 5963 8483
rect 5951 8452 6868 8480
rect 5951 8449 5963 8452
rect 5905 8443 5963 8449
rect 2869 8415 2927 8421
rect 2869 8381 2881 8415
rect 2915 8412 2927 8415
rect 3050 8412 3056 8424
rect 2915 8384 3056 8412
rect 2915 8381 2927 8384
rect 2869 8375 2927 8381
rect 3050 8372 3056 8384
rect 3108 8372 3114 8424
rect 3329 8415 3387 8421
rect 3329 8381 3341 8415
rect 3375 8412 3387 8415
rect 3418 8412 3424 8424
rect 3375 8384 3424 8412
rect 3375 8381 3387 8384
rect 3329 8375 3387 8381
rect 3418 8372 3424 8384
rect 3476 8412 3482 8424
rect 3970 8412 3976 8424
rect 3476 8384 3976 8412
rect 3476 8372 3482 8384
rect 3970 8372 3976 8384
rect 4028 8372 4034 8424
rect 5166 8236 5172 8288
rect 5224 8276 5230 8288
rect 5736 8276 5764 8443
rect 6840 8353 6868 8452
rect 7190 8440 7196 8492
rect 7248 8440 7254 8492
rect 7466 8440 7472 8492
rect 7524 8440 7530 8492
rect 7650 8440 7656 8492
rect 7708 8440 7714 8492
rect 7760 8489 7788 8520
rect 11882 8508 11888 8520
rect 11940 8508 11946 8560
rect 12161 8551 12219 8557
rect 12161 8517 12173 8551
rect 12207 8548 12219 8551
rect 12250 8548 12256 8560
rect 12207 8520 12256 8548
rect 12207 8517 12219 8520
rect 12161 8511 12219 8517
rect 12250 8508 12256 8520
rect 12308 8508 12314 8560
rect 7745 8483 7803 8489
rect 7745 8449 7757 8483
rect 7791 8449 7803 8483
rect 7745 8443 7803 8449
rect 9401 8483 9459 8489
rect 9401 8449 9413 8483
rect 9447 8449 9459 8483
rect 9401 8443 9459 8449
rect 7285 8415 7343 8421
rect 7285 8381 7297 8415
rect 7331 8412 7343 8415
rect 7760 8412 7788 8443
rect 7331 8384 7788 8412
rect 9416 8412 9444 8443
rect 9582 8440 9588 8492
rect 9640 8440 9646 8492
rect 9674 8440 9680 8492
rect 9732 8440 9738 8492
rect 11330 8440 11336 8492
rect 11388 8480 11394 8492
rect 12406 8480 12434 8588
rect 17126 8576 17132 8588
rect 17184 8576 17190 8628
rect 11388 8452 12434 8480
rect 12529 8483 12587 8489
rect 11388 8440 11394 8452
rect 12529 8449 12541 8483
rect 12575 8480 12587 8483
rect 13078 8480 13084 8492
rect 12575 8452 13084 8480
rect 12575 8449 12587 8452
rect 12529 8443 12587 8449
rect 13078 8440 13084 8452
rect 13136 8440 13142 8492
rect 9950 8412 9956 8424
rect 9416 8384 9956 8412
rect 7331 8381 7343 8384
rect 7285 8375 7343 8381
rect 9950 8372 9956 8384
rect 10008 8372 10014 8424
rect 12066 8372 12072 8424
rect 12124 8372 12130 8424
rect 6825 8347 6883 8353
rect 6825 8313 6837 8347
rect 6871 8313 6883 8347
rect 6825 8307 6883 8313
rect 7374 8304 7380 8356
rect 7432 8344 7438 8356
rect 7469 8347 7527 8353
rect 7469 8344 7481 8347
rect 7432 8316 7481 8344
rect 7432 8304 7438 8316
rect 7469 8313 7481 8316
rect 7515 8313 7527 8347
rect 7469 8307 7527 8313
rect 11606 8304 11612 8356
rect 11664 8304 11670 8356
rect 10134 8276 10140 8288
rect 5224 8248 10140 8276
rect 5224 8236 5230 8248
rect 10134 8236 10140 8248
rect 10192 8236 10198 8288
rect 12434 8236 12440 8288
rect 12492 8236 12498 8288
rect 1104 8186 17848 8208
rect 1104 8134 1918 8186
rect 1970 8134 1982 8186
rect 2034 8134 2046 8186
rect 2098 8134 2110 8186
rect 2162 8134 2174 8186
rect 2226 8134 2238 8186
rect 2290 8134 7918 8186
rect 7970 8134 7982 8186
rect 8034 8134 8046 8186
rect 8098 8134 8110 8186
rect 8162 8134 8174 8186
rect 8226 8134 8238 8186
rect 8290 8134 13918 8186
rect 13970 8134 13982 8186
rect 14034 8134 14046 8186
rect 14098 8134 14110 8186
rect 14162 8134 14174 8186
rect 14226 8134 14238 8186
rect 14290 8134 17848 8186
rect 1104 8112 17848 8134
rect 1397 8075 1455 8081
rect 1397 8041 1409 8075
rect 1443 8072 1455 8075
rect 1578 8072 1584 8084
rect 1443 8044 1584 8072
rect 1443 8041 1455 8044
rect 1397 8035 1455 8041
rect 1578 8032 1584 8044
rect 1636 8032 1642 8084
rect 7285 8075 7343 8081
rect 7285 8041 7297 8075
rect 7331 8072 7343 8075
rect 7466 8072 7472 8084
rect 7331 8044 7472 8072
rect 7331 8041 7343 8044
rect 7285 8035 7343 8041
rect 7466 8032 7472 8044
rect 7524 8032 7530 8084
rect 7576 8044 7972 8072
rect 5534 7964 5540 8016
rect 5592 7964 5598 8016
rect 7190 7964 7196 8016
rect 7248 7964 7254 8016
rect 7374 7964 7380 8016
rect 7432 8004 7438 8016
rect 7576 8004 7604 8044
rect 7432 7976 7604 8004
rect 7432 7964 7438 7976
rect 7650 7964 7656 8016
rect 7708 8004 7714 8016
rect 7837 8007 7895 8013
rect 7837 8004 7849 8007
rect 7708 7976 7849 8004
rect 7708 7964 7714 7976
rect 7837 7973 7849 7976
rect 7883 7973 7895 8007
rect 7837 7967 7895 7973
rect 3142 7896 3148 7948
rect 3200 7896 3206 7948
rect 5261 7939 5319 7945
rect 5261 7905 5273 7939
rect 5307 7936 5319 7939
rect 5350 7936 5356 7948
rect 5307 7908 5356 7936
rect 5307 7905 5319 7908
rect 5261 7899 5319 7905
rect 5350 7896 5356 7908
rect 5408 7896 5414 7948
rect 6917 7939 6975 7945
rect 6917 7905 6929 7939
rect 6963 7936 6975 7939
rect 7944 7936 7972 8044
rect 9950 8032 9956 8084
rect 10008 8032 10014 8084
rect 10134 8032 10140 8084
rect 10192 8072 10198 8084
rect 16669 8075 16727 8081
rect 16669 8072 16681 8075
rect 10192 8044 16681 8072
rect 10192 8032 10198 8044
rect 16669 8041 16681 8044
rect 16715 8041 16727 8075
rect 16669 8035 16727 8041
rect 9674 7964 9680 8016
rect 9732 7964 9738 8016
rect 10045 8007 10103 8013
rect 10045 7973 10057 8007
rect 10091 7973 10103 8007
rect 16853 8007 16911 8013
rect 16853 8004 16865 8007
rect 10045 7967 10103 7973
rect 15764 7976 16865 8004
rect 9692 7936 9720 7964
rect 9769 7939 9827 7945
rect 9769 7936 9781 7939
rect 6963 7908 7788 7936
rect 6963 7905 6975 7908
rect 6917 7899 6975 7905
rect 5166 7828 5172 7880
rect 5224 7828 5230 7880
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7868 6883 7871
rect 7374 7868 7380 7880
rect 6871 7840 7380 7868
rect 6871 7837 6883 7840
rect 6825 7831 6883 7837
rect 7374 7828 7380 7840
rect 7432 7828 7438 7880
rect 2314 7760 2320 7812
rect 2372 7760 2378 7812
rect 2869 7803 2927 7809
rect 2869 7769 2881 7803
rect 2915 7800 2927 7803
rect 3418 7800 3424 7812
rect 2915 7772 3424 7800
rect 2915 7769 2927 7772
rect 2869 7763 2927 7769
rect 3418 7760 3424 7772
rect 3476 7760 3482 7812
rect 7760 7809 7788 7908
rect 7852 7908 8248 7936
rect 9692 7908 9781 7936
rect 7852 7880 7880 7908
rect 7834 7828 7840 7880
rect 7892 7828 7898 7880
rect 8220 7877 8248 7908
rect 9769 7905 9781 7908
rect 9815 7905 9827 7939
rect 9769 7899 9827 7905
rect 9950 7896 9956 7948
rect 10008 7936 10014 7948
rect 10060 7936 10088 7967
rect 10008 7908 10088 7936
rect 10008 7896 10014 7908
rect 11054 7896 11060 7948
rect 11112 7896 11118 7948
rect 11333 7939 11391 7945
rect 11333 7905 11345 7939
rect 11379 7936 11391 7939
rect 11790 7936 11796 7948
rect 11379 7908 11796 7936
rect 11379 7905 11391 7908
rect 11333 7899 11391 7905
rect 11790 7896 11796 7908
rect 11848 7896 11854 7948
rect 12066 7896 12072 7948
rect 12124 7936 12130 7948
rect 13081 7939 13139 7945
rect 13081 7936 13093 7939
rect 12124 7908 13093 7936
rect 12124 7896 12130 7908
rect 13081 7905 13093 7908
rect 13127 7905 13139 7939
rect 13081 7899 13139 7905
rect 15764 7880 15792 7976
rect 16853 7973 16865 7976
rect 16899 7973 16911 8007
rect 16853 7967 16911 7973
rect 16761 7939 16819 7945
rect 16761 7936 16773 7939
rect 16500 7908 16773 7936
rect 8112 7871 8170 7877
rect 8112 7837 8124 7871
rect 8158 7837 8170 7871
rect 8112 7831 8170 7837
rect 8205 7871 8263 7877
rect 8205 7837 8217 7871
rect 8251 7837 8263 7871
rect 8205 7831 8263 7837
rect 7745 7803 7803 7809
rect 7745 7769 7757 7803
rect 7791 7769 7803 7803
rect 7745 7763 7803 7769
rect 7760 7732 7788 7763
rect 8128 7732 8156 7831
rect 9490 7828 9496 7880
rect 9548 7868 9554 7880
rect 9677 7871 9735 7877
rect 9677 7868 9689 7871
rect 9548 7840 9689 7868
rect 9548 7828 9554 7840
rect 9677 7837 9689 7840
rect 9723 7837 9735 7871
rect 9677 7831 9735 7837
rect 12434 7828 12440 7880
rect 12492 7828 12498 7880
rect 14458 7828 14464 7880
rect 14516 7868 14522 7880
rect 14829 7871 14887 7877
rect 14829 7868 14841 7871
rect 14516 7840 14841 7868
rect 14516 7828 14522 7840
rect 14829 7837 14841 7840
rect 14875 7837 14887 7871
rect 14829 7831 14887 7837
rect 15746 7828 15752 7880
rect 15804 7828 15810 7880
rect 15930 7877 15936 7880
rect 15903 7871 15936 7877
rect 15903 7837 15915 7871
rect 15903 7831 15936 7837
rect 15930 7828 15936 7831
rect 15988 7828 15994 7880
rect 16500 7877 16528 7908
rect 16761 7905 16773 7908
rect 16807 7905 16819 7939
rect 16761 7899 16819 7905
rect 16117 7871 16175 7877
rect 16117 7837 16129 7871
rect 16163 7868 16175 7871
rect 16209 7871 16267 7877
rect 16209 7868 16221 7871
rect 16163 7840 16221 7868
rect 16163 7837 16175 7840
rect 16117 7831 16175 7837
rect 16209 7837 16221 7840
rect 16255 7837 16267 7871
rect 16209 7831 16267 7837
rect 16485 7871 16543 7877
rect 16485 7837 16497 7871
rect 16531 7837 16543 7871
rect 16485 7831 16543 7837
rect 10134 7760 10140 7812
rect 10192 7800 10198 7812
rect 10413 7803 10471 7809
rect 10413 7800 10425 7803
rect 10192 7772 10425 7800
rect 10192 7760 10198 7772
rect 10413 7769 10425 7772
rect 10459 7769 10471 7803
rect 10413 7763 10471 7769
rect 14366 7760 14372 7812
rect 14424 7800 14430 7812
rect 14645 7803 14703 7809
rect 14645 7800 14657 7803
rect 14424 7772 14657 7800
rect 14424 7760 14430 7772
rect 14645 7769 14657 7772
rect 14691 7769 14703 7803
rect 15948 7800 15976 7828
rect 17221 7803 17279 7809
rect 17221 7800 17233 7803
rect 15948 7772 17233 7800
rect 14645 7763 14703 7769
rect 16500 7744 16528 7772
rect 17221 7769 17233 7772
rect 17267 7769 17279 7803
rect 17221 7763 17279 7769
rect 9309 7735 9367 7741
rect 9309 7732 9321 7735
rect 7760 7704 9321 7732
rect 9309 7701 9321 7704
rect 9355 7701 9367 7735
rect 9309 7695 9367 7701
rect 14461 7735 14519 7741
rect 14461 7701 14473 7735
rect 14507 7732 14519 7735
rect 14550 7732 14556 7744
rect 14507 7704 14556 7732
rect 14507 7701 14519 7704
rect 14461 7695 14519 7701
rect 14550 7692 14556 7704
rect 14608 7692 14614 7744
rect 16206 7692 16212 7744
rect 16264 7732 16270 7744
rect 16301 7735 16359 7741
rect 16301 7732 16313 7735
rect 16264 7704 16313 7732
rect 16264 7692 16270 7704
rect 16301 7701 16313 7704
rect 16347 7701 16359 7735
rect 16301 7695 16359 7701
rect 16482 7692 16488 7744
rect 16540 7692 16546 7744
rect 1104 7642 17848 7664
rect 1104 7590 2658 7642
rect 2710 7590 2722 7642
rect 2774 7590 2786 7642
rect 2838 7590 2850 7642
rect 2902 7590 2914 7642
rect 2966 7590 2978 7642
rect 3030 7590 8658 7642
rect 8710 7590 8722 7642
rect 8774 7590 8786 7642
rect 8838 7590 8850 7642
rect 8902 7590 8914 7642
rect 8966 7590 8978 7642
rect 9030 7590 14658 7642
rect 14710 7590 14722 7642
rect 14774 7590 14786 7642
rect 14838 7590 14850 7642
rect 14902 7590 14914 7642
rect 14966 7590 14978 7642
rect 15030 7590 17848 7642
rect 1104 7568 17848 7590
rect 1302 7488 1308 7540
rect 1360 7528 1366 7540
rect 1397 7531 1455 7537
rect 1397 7528 1409 7531
rect 1360 7500 1409 7528
rect 1360 7488 1366 7500
rect 1397 7497 1409 7500
rect 1443 7497 1455 7531
rect 1397 7491 1455 7497
rect 2314 7488 2320 7540
rect 2372 7488 2378 7540
rect 9490 7488 9496 7540
rect 9548 7488 9554 7540
rect 9582 7488 9588 7540
rect 9640 7488 9646 7540
rect 10134 7488 10140 7540
rect 10192 7488 10198 7540
rect 15565 7531 15623 7537
rect 15565 7497 15577 7531
rect 15611 7528 15623 7531
rect 15746 7528 15752 7540
rect 15611 7500 15752 7528
rect 15611 7497 15623 7500
rect 15565 7491 15623 7497
rect 15746 7488 15752 7500
rect 15804 7488 15810 7540
rect 10152 7460 10180 7488
rect 4448 7432 4936 7460
rect 1578 7352 1584 7404
rect 1636 7352 1642 7404
rect 2406 7352 2412 7404
rect 2464 7352 2470 7404
rect 3789 7395 3847 7401
rect 3789 7361 3801 7395
rect 3835 7392 3847 7395
rect 3878 7392 3884 7404
rect 3835 7364 3884 7392
rect 3835 7361 3847 7364
rect 3789 7355 3847 7361
rect 3878 7352 3884 7364
rect 3936 7392 3942 7404
rect 4448 7401 4476 7432
rect 4433 7395 4491 7401
rect 3936 7364 4108 7392
rect 3936 7352 3942 7364
rect 3418 7284 3424 7336
rect 3476 7284 3482 7336
rect 4080 7333 4108 7364
rect 4433 7361 4445 7395
rect 4479 7361 4491 7395
rect 4709 7395 4767 7401
rect 4709 7392 4721 7395
rect 4433 7355 4491 7361
rect 4540 7364 4721 7392
rect 4540 7333 4568 7364
rect 4709 7361 4721 7364
rect 4755 7392 4767 7395
rect 4798 7392 4804 7404
rect 4755 7364 4804 7392
rect 4755 7361 4767 7364
rect 4709 7355 4767 7361
rect 4798 7352 4804 7364
rect 4856 7352 4862 7404
rect 4908 7401 4936 7432
rect 9140 7432 10180 7460
rect 4893 7395 4951 7401
rect 4893 7361 4905 7395
rect 4939 7392 4951 7395
rect 5810 7392 5816 7404
rect 4939 7364 5816 7392
rect 4939 7361 4951 7364
rect 4893 7355 4951 7361
rect 5810 7352 5816 7364
rect 5868 7352 5874 7404
rect 9140 7401 9168 7432
rect 12434 7420 12440 7472
rect 12492 7420 12498 7472
rect 15102 7420 15108 7472
rect 15160 7460 15166 7472
rect 15160 7432 15240 7460
rect 15160 7420 15166 7432
rect 9125 7395 9183 7401
rect 9125 7361 9137 7395
rect 9171 7361 9183 7395
rect 9125 7355 9183 7361
rect 9766 7352 9772 7404
rect 9824 7352 9830 7404
rect 9950 7352 9956 7404
rect 10008 7352 10014 7404
rect 10045 7395 10103 7401
rect 10045 7361 10057 7395
rect 10091 7361 10103 7395
rect 10045 7355 10103 7361
rect 10229 7395 10287 7401
rect 10229 7361 10241 7395
rect 10275 7392 10287 7395
rect 11054 7392 11060 7404
rect 10275 7364 11060 7392
rect 10275 7361 10287 7364
rect 10229 7355 10287 7361
rect 3697 7327 3755 7333
rect 3697 7293 3709 7327
rect 3743 7293 3755 7327
rect 3697 7287 3755 7293
rect 4065 7327 4123 7333
rect 4065 7293 4077 7327
rect 4111 7293 4123 7327
rect 4065 7287 4123 7293
rect 4525 7327 4583 7333
rect 4525 7293 4537 7327
rect 4571 7293 4583 7327
rect 4525 7287 4583 7293
rect 9217 7327 9275 7333
rect 9217 7293 9229 7327
rect 9263 7293 9275 7327
rect 9784 7324 9812 7352
rect 10060 7324 10088 7355
rect 9784 7296 10088 7324
rect 9217 7287 9275 7293
rect 3712 7256 3740 7287
rect 3786 7256 3792 7268
rect 3712 7228 3792 7256
rect 3786 7216 3792 7228
rect 3844 7216 3850 7268
rect 9232 7256 9260 7287
rect 9858 7256 9864 7268
rect 9232 7228 9864 7256
rect 9858 7216 9864 7228
rect 9916 7216 9922 7268
rect 10244 7256 10272 7355
rect 11054 7352 11060 7364
rect 11112 7352 11118 7404
rect 12158 7352 12164 7404
rect 12216 7352 12222 7404
rect 13538 7352 13544 7404
rect 13596 7352 13602 7404
rect 14366 7352 14372 7404
rect 14424 7392 14430 7404
rect 15212 7401 15240 7432
rect 14553 7395 14611 7401
rect 14553 7392 14565 7395
rect 14424 7364 14565 7392
rect 14424 7352 14430 7364
rect 14553 7361 14565 7364
rect 14599 7361 14611 7395
rect 14553 7355 14611 7361
rect 15197 7395 15255 7401
rect 15197 7361 15209 7395
rect 15243 7361 15255 7395
rect 15197 7355 15255 7361
rect 10873 7327 10931 7333
rect 10873 7293 10885 7327
rect 10919 7324 10931 7327
rect 11238 7324 11244 7336
rect 10919 7296 11244 7324
rect 10919 7293 10931 7296
rect 10873 7287 10931 7293
rect 11238 7284 11244 7296
rect 11296 7324 11302 7336
rect 12066 7324 12072 7336
rect 11296 7296 12072 7324
rect 11296 7284 11302 7296
rect 12066 7284 12072 7296
rect 12124 7284 12130 7336
rect 13630 7284 13636 7336
rect 13688 7324 13694 7336
rect 14185 7327 14243 7333
rect 14185 7324 14197 7327
rect 13688 7296 14197 7324
rect 13688 7284 13694 7296
rect 14185 7293 14197 7296
rect 14231 7293 14243 7327
rect 14185 7287 14243 7293
rect 14458 7284 14464 7336
rect 14516 7324 14522 7336
rect 14642 7324 14648 7336
rect 14516 7296 14648 7324
rect 14516 7284 14522 7296
rect 14642 7284 14648 7296
rect 14700 7284 14706 7336
rect 14921 7327 14979 7333
rect 14921 7293 14933 7327
rect 14967 7324 14979 7327
rect 15105 7327 15163 7333
rect 15105 7324 15117 7327
rect 14967 7296 15117 7324
rect 14967 7293 14979 7296
rect 14921 7287 14979 7293
rect 15105 7293 15117 7296
rect 15151 7293 15163 7327
rect 15764 7324 15792 7488
rect 16482 7352 16488 7404
rect 16540 7392 16546 7404
rect 16853 7395 16911 7401
rect 16853 7392 16865 7395
rect 16540 7364 16865 7392
rect 16540 7352 16546 7364
rect 16853 7361 16865 7364
rect 16899 7361 16911 7395
rect 16853 7355 16911 7361
rect 16761 7327 16819 7333
rect 16761 7324 16773 7327
rect 15764 7296 16773 7324
rect 15105 7287 15163 7293
rect 16761 7293 16773 7296
rect 16807 7293 16819 7327
rect 16761 7287 16819 7293
rect 9968 7228 10272 7256
rect 11149 7259 11207 7265
rect 4706 7148 4712 7200
rect 4764 7148 4770 7200
rect 9968 7197 9996 7228
rect 11149 7225 11161 7259
rect 11195 7256 11207 7259
rect 11422 7256 11428 7268
rect 11195 7228 11428 7256
rect 11195 7225 11207 7228
rect 11149 7219 11207 7225
rect 11422 7216 11428 7228
rect 11480 7216 11486 7268
rect 9953 7191 10011 7197
rect 9953 7157 9965 7191
rect 9999 7157 10011 7191
rect 9953 7151 10011 7157
rect 11333 7191 11391 7197
rect 11333 7157 11345 7191
rect 11379 7188 11391 7191
rect 11514 7188 11520 7200
rect 11379 7160 11520 7188
rect 11379 7157 11391 7160
rect 11333 7151 11391 7157
rect 11514 7148 11520 7160
rect 11572 7148 11578 7200
rect 17218 7148 17224 7200
rect 17276 7148 17282 7200
rect 1104 7098 17848 7120
rect 1104 7046 1918 7098
rect 1970 7046 1982 7098
rect 2034 7046 2046 7098
rect 2098 7046 2110 7098
rect 2162 7046 2174 7098
rect 2226 7046 2238 7098
rect 2290 7046 7918 7098
rect 7970 7046 7982 7098
rect 8034 7046 8046 7098
rect 8098 7046 8110 7098
rect 8162 7046 8174 7098
rect 8226 7046 8238 7098
rect 8290 7046 13918 7098
rect 13970 7046 13982 7098
rect 14034 7046 14046 7098
rect 14098 7046 14110 7098
rect 14162 7046 14174 7098
rect 14226 7046 14238 7098
rect 14290 7046 17848 7098
rect 1104 7024 17848 7046
rect 1397 6987 1455 6993
rect 1397 6953 1409 6987
rect 1443 6984 1455 6987
rect 1578 6984 1584 6996
rect 1443 6956 1584 6984
rect 1443 6953 1455 6956
rect 1397 6947 1455 6953
rect 1578 6944 1584 6956
rect 1636 6944 1642 6996
rect 9950 6944 9956 6996
rect 10008 6984 10014 6996
rect 10594 6984 10600 6996
rect 10008 6956 10600 6984
rect 10008 6944 10014 6956
rect 10594 6944 10600 6956
rect 10652 6944 10658 6996
rect 11054 6944 11060 6996
rect 11112 6944 11118 6996
rect 13725 6987 13783 6993
rect 13725 6953 13737 6987
rect 13771 6984 13783 6987
rect 14366 6984 14372 6996
rect 13771 6956 14372 6984
rect 13771 6953 13783 6956
rect 13725 6947 13783 6953
rect 14366 6944 14372 6956
rect 14424 6984 14430 6996
rect 15194 6984 15200 6996
rect 14424 6956 15200 6984
rect 14424 6944 14430 6956
rect 15194 6944 15200 6956
rect 15252 6944 15258 6996
rect 4798 6876 4804 6928
rect 4856 6916 4862 6928
rect 4856 6888 14964 6916
rect 4856 6876 4862 6888
rect 3142 6808 3148 6860
rect 3200 6808 3206 6860
rect 4154 6808 4160 6860
rect 4212 6848 4218 6860
rect 4249 6851 4307 6857
rect 4249 6848 4261 6851
rect 4212 6820 4261 6848
rect 4212 6808 4218 6820
rect 4249 6817 4261 6820
rect 4295 6817 4307 6851
rect 9122 6848 9128 6860
rect 4249 6811 4307 6817
rect 7392 6820 9128 6848
rect 3786 6740 3792 6792
rect 3844 6740 3850 6792
rect 3878 6740 3884 6792
rect 3936 6740 3942 6792
rect 4065 6783 4123 6789
rect 4065 6749 4077 6783
rect 4111 6780 4123 6783
rect 4706 6780 4712 6792
rect 4111 6752 4712 6780
rect 4111 6749 4123 6752
rect 4065 6743 4123 6749
rect 4706 6740 4712 6752
rect 4764 6740 4770 6792
rect 7392 6789 7420 6820
rect 9122 6808 9128 6820
rect 9180 6808 9186 6860
rect 9309 6851 9367 6857
rect 9309 6817 9321 6851
rect 9355 6848 9367 6851
rect 9766 6848 9772 6860
rect 9355 6820 9772 6848
rect 9355 6817 9367 6820
rect 9309 6811 9367 6817
rect 9766 6808 9772 6820
rect 9824 6808 9830 6860
rect 11422 6808 11428 6860
rect 11480 6848 11486 6860
rect 11701 6851 11759 6857
rect 11480 6820 11652 6848
rect 11480 6808 11486 6820
rect 7377 6783 7435 6789
rect 7377 6749 7389 6783
rect 7423 6749 7435 6783
rect 7377 6743 7435 6749
rect 7466 6740 7472 6792
rect 7524 6780 7530 6792
rect 7653 6783 7711 6789
rect 7653 6780 7665 6783
rect 7524 6752 7665 6780
rect 7524 6740 7530 6752
rect 7653 6749 7665 6752
rect 7699 6749 7711 6783
rect 7653 6743 7711 6749
rect 9217 6783 9275 6789
rect 9217 6749 9229 6783
rect 9263 6749 9275 6783
rect 9217 6743 9275 6749
rect 2314 6672 2320 6724
rect 2372 6672 2378 6724
rect 2869 6715 2927 6721
rect 2869 6681 2881 6715
rect 2915 6712 2927 6715
rect 3602 6712 3608 6724
rect 2915 6684 3608 6712
rect 2915 6681 2927 6684
rect 2869 6675 2927 6681
rect 3602 6672 3608 6684
rect 3660 6672 3666 6724
rect 7558 6672 7564 6724
rect 7616 6672 7622 6724
rect 8570 6604 8576 6656
rect 8628 6644 8634 6656
rect 9238 6644 9266 6743
rect 9398 6740 9404 6792
rect 9456 6740 9462 6792
rect 11440 6780 11468 6808
rect 9508 6752 11468 6780
rect 9306 6672 9312 6724
rect 9364 6712 9370 6724
rect 9508 6712 9536 6752
rect 11514 6740 11520 6792
rect 11572 6740 11578 6792
rect 11624 6780 11652 6820
rect 11701 6817 11713 6851
rect 11747 6848 11759 6851
rect 12250 6848 12256 6860
rect 11747 6820 12256 6848
rect 11747 6817 11759 6820
rect 11701 6811 11759 6817
rect 12250 6808 12256 6820
rect 12308 6848 12314 6860
rect 12618 6848 12624 6860
rect 12308 6820 12624 6848
rect 12308 6808 12314 6820
rect 12618 6808 12624 6820
rect 12676 6808 12682 6860
rect 13357 6851 13415 6857
rect 13357 6817 13369 6851
rect 13403 6848 13415 6851
rect 13538 6848 13544 6860
rect 13403 6820 13544 6848
rect 13403 6817 13415 6820
rect 13357 6811 13415 6817
rect 13538 6808 13544 6820
rect 13596 6808 13602 6860
rect 13633 6851 13691 6857
rect 13633 6817 13645 6851
rect 13679 6817 13691 6851
rect 13633 6811 13691 6817
rect 11885 6783 11943 6789
rect 11885 6780 11897 6783
rect 11624 6752 11897 6780
rect 11885 6749 11897 6752
rect 11931 6749 11943 6783
rect 11885 6743 11943 6749
rect 12066 6740 12072 6792
rect 12124 6740 12130 6792
rect 12158 6740 12164 6792
rect 12216 6780 12222 6792
rect 12216 6752 12434 6780
rect 12216 6740 12222 6752
rect 9364 6684 9536 6712
rect 11425 6715 11483 6721
rect 9364 6672 9370 6684
rect 11425 6681 11437 6715
rect 11471 6712 11483 6715
rect 11606 6712 11612 6724
rect 11471 6684 11612 6712
rect 11471 6681 11483 6684
rect 11425 6675 11483 6681
rect 11606 6672 11612 6684
rect 11664 6712 11670 6724
rect 12253 6715 12311 6721
rect 12253 6712 12265 6715
rect 11664 6684 12265 6712
rect 11664 6672 11670 6684
rect 12253 6681 12265 6684
rect 12299 6681 12311 6715
rect 12406 6712 12434 6752
rect 13078 6740 13084 6792
rect 13136 6780 13142 6792
rect 13449 6783 13507 6789
rect 13449 6780 13461 6783
rect 13136 6752 13461 6780
rect 13136 6740 13142 6752
rect 13449 6749 13461 6752
rect 13495 6749 13507 6783
rect 13449 6743 13507 6749
rect 13648 6712 13676 6811
rect 14366 6808 14372 6860
rect 14424 6808 14430 6860
rect 14936 6848 14964 6888
rect 16393 6851 16451 6857
rect 16393 6848 16405 6851
rect 14936 6820 16405 6848
rect 16393 6817 16405 6820
rect 16439 6817 16451 6851
rect 16393 6811 16451 6817
rect 17218 6808 17224 6860
rect 17276 6808 17282 6860
rect 13814 6740 13820 6792
rect 13872 6740 13878 6792
rect 13909 6783 13967 6789
rect 13909 6749 13921 6783
rect 13955 6780 13967 6783
rect 13998 6780 14004 6792
rect 13955 6752 14004 6780
rect 13955 6749 13967 6752
rect 13909 6743 13967 6749
rect 13998 6740 14004 6752
rect 14056 6740 14062 6792
rect 14550 6740 14556 6792
rect 14608 6740 14614 6792
rect 14734 6740 14740 6792
rect 14792 6740 14798 6792
rect 14829 6783 14887 6789
rect 14829 6749 14841 6783
rect 14875 6780 14887 6783
rect 15010 6780 15016 6792
rect 14875 6752 15016 6780
rect 14875 6749 14887 6752
rect 14829 6743 14887 6749
rect 15010 6740 15016 6752
rect 15068 6740 15074 6792
rect 15105 6783 15163 6789
rect 15105 6749 15117 6783
rect 15151 6749 15163 6783
rect 15105 6743 15163 6749
rect 12406 6684 13676 6712
rect 12253 6675 12311 6681
rect 14642 6672 14648 6724
rect 14700 6712 14706 6724
rect 15120 6712 15148 6743
rect 15194 6740 15200 6792
rect 15252 6740 15258 6792
rect 16206 6740 16212 6792
rect 16264 6780 16270 6792
rect 17037 6783 17095 6789
rect 17037 6780 17049 6783
rect 16264 6752 17049 6780
rect 16264 6740 16270 6752
rect 17037 6749 17049 6752
rect 17083 6749 17095 6783
rect 17037 6743 17095 6749
rect 14700 6684 15148 6712
rect 14700 6672 14706 6684
rect 15120 6656 15148 6684
rect 13906 6644 13912 6656
rect 8628 6616 13912 6644
rect 8628 6604 8634 6616
rect 13906 6604 13912 6616
rect 13964 6644 13970 6656
rect 14366 6644 14372 6656
rect 13964 6616 14372 6644
rect 13964 6604 13970 6616
rect 14366 6604 14372 6616
rect 14424 6604 14430 6656
rect 14734 6604 14740 6656
rect 14792 6644 14798 6656
rect 14921 6647 14979 6653
rect 14921 6644 14933 6647
rect 14792 6616 14933 6644
rect 14792 6604 14798 6616
rect 14921 6613 14933 6616
rect 14967 6613 14979 6647
rect 14921 6607 14979 6613
rect 15102 6604 15108 6656
rect 15160 6604 15166 6656
rect 1104 6554 17848 6576
rect 1104 6502 2658 6554
rect 2710 6502 2722 6554
rect 2774 6502 2786 6554
rect 2838 6502 2850 6554
rect 2902 6502 2914 6554
rect 2966 6502 2978 6554
rect 3030 6502 8658 6554
rect 8710 6502 8722 6554
rect 8774 6502 8786 6554
rect 8838 6502 8850 6554
rect 8902 6502 8914 6554
rect 8966 6502 8978 6554
rect 9030 6502 14658 6554
rect 14710 6502 14722 6554
rect 14774 6502 14786 6554
rect 14838 6502 14850 6554
rect 14902 6502 14914 6554
rect 14966 6502 14978 6554
rect 15030 6502 17848 6554
rect 1104 6480 17848 6502
rect 1302 6400 1308 6452
rect 1360 6440 1366 6452
rect 1397 6443 1455 6449
rect 1397 6440 1409 6443
rect 1360 6412 1409 6440
rect 1360 6400 1366 6412
rect 1397 6409 1409 6412
rect 1443 6409 1455 6443
rect 1397 6403 1455 6409
rect 2314 6400 2320 6452
rect 2372 6400 2378 6452
rect 3786 6400 3792 6452
rect 3844 6440 3850 6452
rect 4709 6443 4767 6449
rect 4709 6440 4721 6443
rect 3844 6412 4721 6440
rect 3844 6400 3850 6412
rect 4709 6409 4721 6412
rect 4755 6409 4767 6443
rect 4709 6403 4767 6409
rect 5810 6400 5816 6452
rect 5868 6400 5874 6452
rect 9125 6443 9183 6449
rect 9125 6409 9137 6443
rect 9171 6409 9183 6443
rect 9125 6403 9183 6409
rect 3988 6344 4384 6372
rect 1578 6264 1584 6316
rect 1636 6264 1642 6316
rect 2406 6264 2412 6316
rect 2464 6264 2470 6316
rect 3988 6313 4016 6344
rect 4356 6316 4384 6344
rect 7650 6332 7656 6384
rect 7708 6372 7714 6384
rect 8665 6375 8723 6381
rect 8665 6372 8677 6375
rect 7708 6344 8677 6372
rect 7708 6332 7714 6344
rect 8665 6341 8677 6344
rect 8711 6341 8723 6375
rect 9140 6372 9168 6403
rect 10134 6400 10140 6452
rect 10192 6440 10198 6452
rect 16298 6440 16304 6452
rect 10192 6412 16304 6440
rect 10192 6400 10198 6412
rect 16298 6400 16304 6412
rect 16356 6400 16362 6452
rect 11882 6372 11888 6384
rect 9140 6344 11888 6372
rect 8665 6335 8723 6341
rect 11882 6332 11888 6344
rect 11940 6332 11946 6384
rect 12250 6332 12256 6384
rect 12308 6372 12314 6384
rect 12713 6375 12771 6381
rect 12713 6372 12725 6375
rect 12308 6344 12725 6372
rect 12308 6332 12314 6344
rect 12713 6341 12725 6344
rect 12759 6372 12771 6375
rect 14274 6372 14280 6384
rect 12759 6344 14280 6372
rect 12759 6341 12771 6344
rect 12713 6335 12771 6341
rect 14274 6332 14280 6344
rect 14332 6332 14338 6384
rect 14366 6332 14372 6384
rect 14424 6372 14430 6384
rect 14424 6344 14780 6372
rect 14424 6332 14430 6344
rect 3973 6307 4031 6313
rect 3973 6273 3985 6307
rect 4019 6273 4031 6307
rect 4246 6304 4252 6316
rect 3973 6267 4031 6273
rect 4080 6276 4252 6304
rect 3602 6196 3608 6248
rect 3660 6196 3666 6248
rect 4080 6245 4108 6276
rect 4246 6264 4252 6276
rect 4304 6264 4310 6316
rect 4338 6264 4344 6316
rect 4396 6264 4402 6316
rect 4525 6307 4583 6313
rect 4525 6273 4537 6307
rect 4571 6304 4583 6307
rect 5902 6304 5908 6316
rect 4571 6276 5908 6304
rect 4571 6273 4583 6276
rect 4525 6267 4583 6273
rect 5902 6264 5908 6276
rect 5960 6264 5966 6316
rect 6088 6307 6146 6313
rect 6088 6273 6100 6307
rect 6134 6273 6146 6307
rect 6088 6267 6146 6273
rect 6181 6307 6239 6313
rect 6181 6273 6193 6307
rect 6227 6304 6239 6307
rect 6730 6304 6736 6316
rect 6227 6276 6736 6304
rect 6227 6273 6239 6276
rect 6181 6267 6239 6273
rect 4065 6239 4123 6245
rect 4065 6205 4077 6239
rect 4111 6205 4123 6239
rect 6104 6236 6132 6267
rect 6730 6264 6736 6276
rect 6788 6264 6794 6316
rect 7374 6264 7380 6316
rect 7432 6304 7438 6316
rect 7929 6307 7987 6313
rect 7929 6304 7941 6307
rect 7432 6276 7941 6304
rect 7432 6264 7438 6276
rect 7929 6273 7941 6276
rect 7975 6273 7987 6307
rect 7929 6267 7987 6273
rect 8113 6307 8171 6313
rect 8113 6273 8125 6307
rect 8159 6273 8171 6307
rect 8113 6267 8171 6273
rect 6825 6239 6883 6245
rect 6825 6236 6837 6239
rect 6104 6208 6837 6236
rect 4065 6199 4123 6205
rect 6825 6205 6837 6208
rect 6871 6236 6883 6239
rect 7742 6236 7748 6248
rect 6871 6208 7748 6236
rect 6871 6205 6883 6208
rect 6825 6199 6883 6205
rect 7742 6196 7748 6208
rect 7800 6196 7806 6248
rect 8128 6168 8156 6267
rect 8386 6264 8392 6316
rect 8444 6304 8450 6316
rect 8757 6307 8815 6313
rect 8757 6304 8769 6307
rect 8444 6276 8769 6304
rect 8444 6264 8450 6276
rect 8757 6273 8769 6276
rect 8803 6273 8815 6307
rect 8757 6267 8815 6273
rect 9858 6264 9864 6316
rect 9916 6264 9922 6316
rect 11606 6264 11612 6316
rect 11664 6304 11670 6316
rect 11977 6307 12035 6313
rect 11977 6304 11989 6307
rect 11664 6276 11989 6304
rect 11664 6264 11670 6276
rect 11977 6273 11989 6276
rect 12023 6273 12035 6307
rect 11977 6267 12035 6273
rect 12618 6264 12624 6316
rect 12676 6304 12682 6316
rect 12897 6307 12955 6313
rect 12676 6276 12721 6304
rect 12676 6264 12682 6276
rect 12897 6273 12909 6307
rect 12943 6304 12955 6307
rect 14461 6307 14519 6313
rect 14461 6304 14473 6307
rect 12943 6276 14473 6304
rect 12943 6273 12955 6276
rect 12897 6267 12955 6273
rect 14461 6273 14473 6276
rect 14507 6273 14519 6307
rect 14461 6267 14519 6273
rect 8570 6196 8576 6248
rect 8628 6196 8634 6248
rect 10134 6196 10140 6248
rect 10192 6196 10198 6248
rect 11790 6196 11796 6248
rect 11848 6196 11854 6248
rect 11885 6239 11943 6245
rect 11885 6205 11897 6239
rect 11931 6205 11943 6239
rect 11885 6199 11943 6205
rect 11514 6168 11520 6180
rect 8128 6140 11520 6168
rect 11514 6128 11520 6140
rect 11572 6168 11578 6180
rect 11900 6168 11928 6199
rect 12434 6196 12440 6248
rect 12492 6236 12498 6248
rect 12912 6236 12940 6267
rect 14550 6264 14556 6316
rect 14608 6304 14614 6316
rect 14752 6313 14780 6344
rect 14645 6307 14703 6313
rect 14645 6304 14657 6307
rect 14608 6276 14657 6304
rect 14608 6264 14614 6276
rect 14645 6273 14657 6276
rect 14691 6273 14703 6307
rect 14645 6267 14703 6273
rect 14737 6307 14795 6313
rect 14737 6273 14749 6307
rect 14783 6304 14795 6307
rect 14826 6304 14832 6316
rect 14783 6276 14832 6304
rect 14783 6273 14795 6276
rect 14737 6267 14795 6273
rect 14826 6264 14832 6276
rect 14884 6264 14890 6316
rect 12492 6208 12940 6236
rect 12492 6196 12498 6208
rect 11572 6140 11928 6168
rect 12345 6171 12403 6177
rect 11572 6128 11578 6140
rect 12345 6137 12357 6171
rect 12391 6168 12403 6171
rect 15930 6168 15936 6180
rect 12391 6140 15936 6168
rect 12391 6137 12403 6140
rect 12345 6131 12403 6137
rect 15930 6128 15936 6140
rect 15988 6128 15994 6180
rect 6362 6060 6368 6112
rect 6420 6100 6426 6112
rect 6457 6103 6515 6109
rect 6457 6100 6469 6103
rect 6420 6072 6469 6100
rect 6420 6060 6426 6072
rect 6457 6069 6469 6072
rect 6503 6069 6515 6103
rect 6457 6063 6515 6069
rect 7834 6060 7840 6112
rect 7892 6100 7898 6112
rect 8021 6103 8079 6109
rect 8021 6100 8033 6103
rect 7892 6072 8033 6100
rect 7892 6060 7898 6072
rect 8021 6069 8033 6072
rect 8067 6069 8079 6103
rect 8021 6063 8079 6069
rect 9950 6060 9956 6112
rect 10008 6060 10014 6112
rect 10042 6060 10048 6112
rect 10100 6060 10106 6112
rect 11882 6060 11888 6112
rect 11940 6100 11946 6112
rect 12618 6100 12624 6112
rect 11940 6072 12624 6100
rect 11940 6060 11946 6072
rect 12618 6060 12624 6072
rect 12676 6060 12682 6112
rect 12802 6060 12808 6112
rect 12860 6100 12866 6112
rect 12897 6103 12955 6109
rect 12897 6100 12909 6103
rect 12860 6072 12909 6100
rect 12860 6060 12866 6072
rect 12897 6069 12909 6072
rect 12943 6069 12955 6103
rect 12897 6063 12955 6069
rect 14366 6060 14372 6112
rect 14424 6100 14430 6112
rect 14461 6103 14519 6109
rect 14461 6100 14473 6103
rect 14424 6072 14473 6100
rect 14424 6060 14430 6072
rect 14461 6069 14473 6072
rect 14507 6069 14519 6103
rect 14461 6063 14519 6069
rect 1104 6010 17848 6032
rect 1104 5958 1918 6010
rect 1970 5958 1982 6010
rect 2034 5958 2046 6010
rect 2098 5958 2110 6010
rect 2162 5958 2174 6010
rect 2226 5958 2238 6010
rect 2290 5958 7918 6010
rect 7970 5958 7982 6010
rect 8034 5958 8046 6010
rect 8098 5958 8110 6010
rect 8162 5958 8174 6010
rect 8226 5958 8238 6010
rect 8290 5958 13918 6010
rect 13970 5958 13982 6010
rect 14034 5958 14046 6010
rect 14098 5958 14110 6010
rect 14162 5958 14174 6010
rect 14226 5958 14238 6010
rect 14290 5958 17848 6010
rect 1104 5936 17848 5958
rect 4246 5856 4252 5908
rect 4304 5856 4310 5908
rect 4338 5856 4344 5908
rect 4396 5896 4402 5908
rect 5629 5899 5687 5905
rect 5629 5896 5641 5899
rect 4396 5868 5641 5896
rect 4396 5856 4402 5868
rect 5629 5865 5641 5868
rect 5675 5865 5687 5899
rect 5629 5859 5687 5865
rect 5902 5856 5908 5908
rect 5960 5896 5966 5908
rect 6181 5899 6239 5905
rect 6181 5896 6193 5899
rect 5960 5868 6193 5896
rect 5960 5856 5966 5868
rect 6181 5865 6193 5868
rect 6227 5865 6239 5899
rect 6181 5859 6239 5865
rect 7650 5856 7656 5908
rect 7708 5856 7714 5908
rect 7742 5856 7748 5908
rect 7800 5896 7806 5908
rect 9585 5899 9643 5905
rect 9585 5896 9597 5899
rect 7800 5868 9597 5896
rect 7800 5856 7806 5868
rect 9585 5865 9597 5868
rect 9631 5865 9643 5899
rect 9585 5859 9643 5865
rect 9950 5856 9956 5908
rect 10008 5896 10014 5908
rect 10321 5899 10379 5905
rect 10321 5896 10333 5899
rect 10008 5868 10333 5896
rect 10008 5856 10014 5868
rect 10321 5865 10333 5868
rect 10367 5896 10379 5899
rect 10410 5896 10416 5908
rect 10367 5868 10416 5896
rect 10367 5865 10379 5868
rect 10321 5859 10379 5865
rect 10410 5856 10416 5868
rect 10468 5856 10474 5908
rect 10505 5899 10563 5905
rect 10505 5865 10517 5899
rect 10551 5865 10563 5899
rect 10505 5859 10563 5865
rect 6362 5828 6368 5840
rect 6012 5800 6368 5828
rect 6012 5769 6040 5800
rect 6362 5788 6368 5800
rect 6420 5788 6426 5840
rect 7098 5788 7104 5840
rect 7156 5828 7162 5840
rect 8202 5828 8208 5840
rect 7156 5800 8208 5828
rect 7156 5788 7162 5800
rect 8202 5788 8208 5800
rect 8260 5788 8266 5840
rect 9214 5788 9220 5840
rect 9272 5788 9278 5840
rect 9493 5831 9551 5837
rect 9493 5797 9505 5831
rect 9539 5828 9551 5831
rect 9858 5828 9864 5840
rect 9539 5800 9864 5828
rect 9539 5797 9551 5800
rect 9493 5791 9551 5797
rect 9858 5788 9864 5800
rect 9916 5828 9922 5840
rect 10226 5828 10232 5840
rect 9916 5800 10232 5828
rect 9916 5788 9922 5800
rect 10226 5788 10232 5800
rect 10284 5788 10290 5840
rect 10520 5828 10548 5859
rect 11146 5856 11152 5908
rect 11204 5856 11210 5908
rect 12437 5899 12495 5905
rect 12437 5896 12449 5899
rect 11256 5868 12449 5896
rect 10336 5800 10548 5828
rect 5997 5763 6055 5769
rect 5997 5729 6009 5763
rect 6043 5729 6055 5763
rect 5997 5723 6055 5729
rect 7374 5720 7380 5772
rect 7432 5760 7438 5772
rect 9232 5760 9260 5788
rect 10336 5772 10364 5800
rect 10594 5788 10600 5840
rect 10652 5828 10658 5840
rect 11256 5828 11284 5868
rect 12437 5865 12449 5868
rect 12483 5865 12495 5899
rect 12437 5859 12495 5865
rect 12618 5856 12624 5908
rect 12676 5896 12682 5908
rect 13081 5899 13139 5905
rect 13081 5896 13093 5899
rect 12676 5868 13093 5896
rect 12676 5856 12682 5868
rect 13081 5865 13093 5868
rect 13127 5865 13139 5899
rect 13081 5859 13139 5865
rect 16206 5856 16212 5908
rect 16264 5856 16270 5908
rect 16482 5856 16488 5908
rect 16540 5856 16546 5908
rect 12158 5828 12164 5840
rect 10652 5800 11284 5828
rect 11624 5800 12164 5828
rect 10652 5788 10658 5800
rect 10318 5760 10324 5772
rect 7432 5732 9260 5760
rect 9324 5732 10324 5760
rect 7432 5720 7438 5732
rect 1486 5652 1492 5704
rect 1544 5692 1550 5704
rect 1581 5695 1639 5701
rect 1581 5692 1593 5695
rect 1544 5664 1593 5692
rect 1544 5652 1550 5664
rect 1581 5661 1593 5664
rect 1627 5661 1639 5695
rect 1581 5655 1639 5661
rect 4430 5652 4436 5704
rect 4488 5652 4494 5704
rect 4614 5652 4620 5704
rect 4672 5692 4678 5704
rect 4709 5695 4767 5701
rect 4709 5692 4721 5695
rect 4672 5664 4721 5692
rect 4672 5652 4678 5664
rect 4709 5661 4721 5664
rect 4755 5661 4767 5695
rect 4709 5655 4767 5661
rect 5905 5695 5963 5701
rect 5905 5661 5917 5695
rect 5951 5661 5963 5695
rect 5905 5655 5963 5661
rect 5920 5624 5948 5655
rect 7466 5652 7472 5704
rect 7524 5652 7530 5704
rect 7623 5695 7681 5701
rect 7623 5661 7635 5695
rect 7669 5692 7681 5695
rect 7669 5664 7880 5692
rect 7669 5661 7681 5664
rect 7623 5655 7681 5661
rect 6638 5624 6644 5636
rect 5920 5596 6644 5624
rect 6638 5584 6644 5596
rect 6696 5584 6702 5636
rect 7852 5624 7880 5664
rect 7926 5652 7932 5704
rect 7984 5652 7990 5704
rect 8110 5652 8116 5704
rect 8168 5652 8174 5704
rect 8202 5652 8208 5704
rect 8260 5652 8266 5704
rect 8294 5652 8300 5704
rect 8352 5652 8358 5704
rect 8496 5701 8524 5732
rect 9324 5701 9352 5732
rect 10318 5720 10324 5732
rect 10376 5720 10382 5772
rect 11624 5769 11652 5800
rect 12158 5788 12164 5800
rect 12216 5828 12222 5840
rect 12216 5800 13584 5828
rect 12216 5788 12222 5800
rect 11609 5763 11667 5769
rect 11609 5729 11621 5763
rect 11655 5729 11667 5763
rect 11609 5723 11667 5729
rect 11701 5763 11759 5769
rect 11701 5729 11713 5763
rect 11747 5760 11759 5763
rect 11882 5760 11888 5772
rect 11747 5732 11888 5760
rect 11747 5729 11759 5732
rect 11701 5723 11759 5729
rect 11882 5720 11888 5732
rect 11940 5720 11946 5772
rect 12272 5763 12330 5769
rect 12272 5729 12284 5763
rect 12318 5760 12330 5763
rect 12318 5732 12756 5760
rect 12318 5729 12330 5732
rect 12272 5723 12330 5729
rect 8481 5695 8539 5701
rect 8481 5661 8493 5695
rect 8527 5661 8539 5695
rect 8481 5655 8539 5661
rect 9217 5695 9275 5701
rect 9217 5661 9229 5695
rect 9263 5661 9275 5695
rect 9217 5655 9275 5661
rect 9309 5695 9367 5701
rect 9309 5661 9321 5695
rect 9355 5661 9367 5695
rect 9309 5655 9367 5661
rect 9122 5624 9128 5636
rect 7852 5596 9128 5624
rect 9122 5584 9128 5596
rect 9180 5584 9186 5636
rect 1394 5516 1400 5568
rect 1452 5516 1458 5568
rect 4154 5516 4160 5568
rect 4212 5556 4218 5568
rect 4617 5559 4675 5565
rect 4617 5556 4629 5559
rect 4212 5528 4629 5556
rect 4212 5516 4218 5528
rect 4617 5525 4629 5528
rect 4663 5525 4675 5559
rect 4617 5519 4675 5525
rect 7190 5516 7196 5568
rect 7248 5556 7254 5568
rect 7558 5556 7564 5568
rect 7248 5528 7564 5556
rect 7248 5516 7254 5528
rect 7558 5516 7564 5528
rect 7616 5556 7622 5568
rect 8110 5556 8116 5568
rect 7616 5528 8116 5556
rect 7616 5516 7622 5528
rect 8110 5516 8116 5528
rect 8168 5516 8174 5568
rect 8478 5516 8484 5568
rect 8536 5556 8542 5568
rect 8665 5559 8723 5565
rect 8665 5556 8677 5559
rect 8536 5528 8677 5556
rect 8536 5516 8542 5528
rect 8665 5525 8677 5528
rect 8711 5525 8723 5559
rect 9232 5556 9260 5655
rect 9766 5652 9772 5704
rect 9824 5652 9830 5704
rect 9861 5695 9919 5701
rect 9861 5661 9873 5695
rect 9907 5692 9919 5695
rect 9907 5664 10732 5692
rect 9907 5661 9919 5664
rect 9861 5655 9919 5661
rect 9493 5627 9551 5633
rect 9493 5593 9505 5627
rect 9539 5624 9551 5627
rect 9876 5624 9904 5655
rect 10704 5636 10732 5664
rect 11790 5652 11796 5704
rect 11848 5692 11854 5704
rect 12069 5695 12127 5701
rect 12069 5692 12081 5695
rect 11848 5664 12081 5692
rect 11848 5652 11854 5664
rect 12069 5661 12081 5664
rect 12115 5692 12127 5695
rect 12115 5664 12572 5692
rect 12115 5661 12127 5664
rect 12069 5655 12127 5661
rect 9539 5596 9904 5624
rect 9968 5596 10456 5624
rect 9539 5593 9551 5596
rect 9493 5587 9551 5593
rect 9766 5556 9772 5568
rect 9232 5528 9772 5556
rect 8665 5519 8723 5525
rect 9766 5516 9772 5528
rect 9824 5556 9830 5568
rect 9968 5556 9996 5596
rect 9824 5528 9996 5556
rect 10229 5559 10287 5565
rect 9824 5516 9830 5528
rect 10229 5525 10241 5559
rect 10275 5556 10287 5559
rect 10318 5556 10324 5568
rect 10275 5528 10324 5556
rect 10275 5525 10287 5528
rect 10229 5519 10287 5525
rect 10318 5516 10324 5528
rect 10376 5516 10382 5568
rect 10428 5556 10456 5596
rect 10686 5584 10692 5636
rect 10744 5584 10750 5636
rect 12161 5627 12219 5633
rect 12161 5593 12173 5627
rect 12207 5624 12219 5627
rect 12250 5624 12256 5636
rect 12207 5596 12256 5624
rect 12207 5593 12219 5596
rect 12161 5587 12219 5593
rect 12250 5584 12256 5596
rect 12308 5584 12314 5636
rect 12342 5584 12348 5636
rect 12400 5584 12406 5636
rect 12544 5624 12572 5664
rect 12618 5652 12624 5704
rect 12676 5652 12682 5704
rect 12728 5701 12756 5732
rect 12894 5720 12900 5772
rect 12952 5720 12958 5772
rect 13446 5760 13452 5772
rect 13004 5732 13452 5760
rect 13004 5701 13032 5732
rect 13446 5720 13452 5732
rect 13504 5720 13510 5772
rect 13556 5769 13584 5800
rect 14274 5788 14280 5840
rect 14332 5828 14338 5840
rect 14921 5831 14979 5837
rect 14921 5828 14933 5831
rect 14332 5800 14933 5828
rect 14332 5788 14338 5800
rect 14921 5797 14933 5800
rect 14967 5797 14979 5831
rect 16574 5828 16580 5840
rect 14921 5791 14979 5797
rect 15948 5800 16580 5828
rect 13541 5763 13599 5769
rect 13541 5729 13553 5763
rect 13587 5729 13599 5763
rect 13541 5723 13599 5729
rect 12713 5695 12771 5701
rect 12713 5661 12725 5695
rect 12759 5661 12771 5695
rect 12713 5655 12771 5661
rect 12989 5695 13047 5701
rect 12989 5661 13001 5695
rect 13035 5661 13047 5695
rect 13556 5692 13584 5723
rect 13722 5720 13728 5772
rect 13780 5720 13786 5772
rect 14642 5720 14648 5772
rect 14700 5760 14706 5772
rect 14737 5763 14795 5769
rect 14737 5760 14749 5763
rect 14700 5732 14749 5760
rect 14700 5720 14706 5732
rect 14737 5729 14749 5732
rect 14783 5760 14795 5763
rect 14826 5760 14832 5772
rect 14783 5732 14832 5760
rect 14783 5729 14795 5732
rect 14737 5723 14795 5729
rect 14826 5720 14832 5732
rect 14884 5720 14890 5772
rect 15562 5720 15568 5772
rect 15620 5720 15626 5772
rect 14553 5695 14611 5701
rect 14553 5692 14565 5695
rect 13556 5664 14565 5692
rect 12989 5655 13047 5661
rect 14553 5661 14565 5664
rect 14599 5692 14611 5695
rect 15378 5692 15384 5704
rect 14599 5664 15384 5692
rect 14599 5661 14611 5664
rect 14553 5655 14611 5661
rect 13004 5624 13032 5655
rect 15378 5652 15384 5664
rect 15436 5652 15442 5704
rect 15948 5701 15976 5800
rect 16574 5788 16580 5800
rect 16632 5788 16638 5840
rect 16117 5763 16175 5769
rect 16117 5729 16129 5763
rect 16163 5760 16175 5763
rect 16390 5760 16396 5772
rect 16163 5732 16396 5760
rect 16163 5729 16175 5732
rect 16117 5723 16175 5729
rect 16390 5720 16396 5732
rect 16448 5720 16454 5772
rect 16666 5720 16672 5772
rect 16724 5720 16730 5772
rect 15933 5695 15991 5701
rect 15933 5661 15945 5695
rect 15979 5661 15991 5695
rect 16408 5692 16436 5720
rect 16761 5695 16819 5701
rect 16761 5692 16773 5695
rect 16408 5664 16773 5692
rect 15933 5655 15991 5661
rect 16761 5661 16773 5664
rect 16807 5661 16819 5695
rect 16761 5655 16819 5661
rect 12544 5596 13032 5624
rect 13446 5584 13452 5636
rect 13504 5624 13510 5636
rect 14461 5627 14519 5633
rect 14461 5624 14473 5627
rect 13504 5596 14473 5624
rect 13504 5584 13510 5596
rect 14461 5593 14473 5596
rect 14507 5624 14519 5627
rect 15289 5627 15347 5633
rect 15289 5624 15301 5627
rect 14507 5596 15301 5624
rect 14507 5593 14519 5596
rect 14461 5587 14519 5593
rect 15289 5593 15301 5596
rect 15335 5593 15347 5627
rect 15289 5587 15347 5593
rect 16298 5584 16304 5636
rect 16356 5584 16362 5636
rect 10489 5559 10547 5565
rect 10489 5556 10501 5559
rect 10428 5528 10501 5556
rect 10489 5525 10501 5528
rect 10535 5556 10547 5559
rect 10870 5556 10876 5568
rect 10535 5528 10876 5556
rect 10535 5525 10547 5528
rect 10489 5519 10547 5525
rect 10870 5516 10876 5528
rect 10928 5516 10934 5568
rect 11054 5516 11060 5568
rect 11112 5556 11118 5568
rect 11517 5559 11575 5565
rect 11517 5556 11529 5559
rect 11112 5528 11529 5556
rect 11112 5516 11118 5528
rect 11517 5525 11529 5528
rect 11563 5525 11575 5559
rect 11517 5519 11575 5525
rect 14090 5516 14096 5568
rect 14148 5516 14154 5568
rect 1104 5466 17848 5488
rect 1104 5414 2658 5466
rect 2710 5414 2722 5466
rect 2774 5414 2786 5466
rect 2838 5414 2850 5466
rect 2902 5414 2914 5466
rect 2966 5414 2978 5466
rect 3030 5414 8658 5466
rect 8710 5414 8722 5466
rect 8774 5414 8786 5466
rect 8838 5414 8850 5466
rect 8902 5414 8914 5466
rect 8966 5414 8978 5466
rect 9030 5414 14658 5466
rect 14710 5414 14722 5466
rect 14774 5414 14786 5466
rect 14838 5414 14850 5466
rect 14902 5414 14914 5466
rect 14966 5414 14978 5466
rect 15030 5414 17848 5466
rect 1104 5392 17848 5414
rect 1397 5355 1455 5361
rect 1397 5321 1409 5355
rect 1443 5352 1455 5355
rect 1578 5352 1584 5364
rect 1443 5324 1584 5352
rect 1443 5321 1455 5324
rect 1397 5315 1455 5321
rect 1578 5312 1584 5324
rect 1636 5312 1642 5364
rect 5353 5355 5411 5361
rect 5353 5321 5365 5355
rect 5399 5352 5411 5355
rect 5810 5352 5816 5364
rect 5399 5324 5816 5352
rect 5399 5321 5411 5324
rect 5353 5315 5411 5321
rect 5810 5312 5816 5324
rect 5868 5312 5874 5364
rect 7745 5355 7803 5361
rect 7745 5321 7757 5355
rect 7791 5321 7803 5355
rect 7745 5315 7803 5321
rect 8113 5355 8171 5361
rect 8113 5321 8125 5355
rect 8159 5352 8171 5355
rect 8294 5352 8300 5364
rect 8159 5324 8300 5352
rect 8159 5321 8171 5324
rect 8113 5315 8171 5321
rect 2314 5244 2320 5296
rect 2372 5244 2378 5296
rect 4430 5244 4436 5296
rect 4488 5284 4494 5296
rect 5689 5287 5747 5293
rect 5689 5284 5701 5287
rect 4488 5256 4752 5284
rect 4488 5244 4494 5256
rect 3142 5176 3148 5228
rect 3200 5176 3206 5228
rect 3881 5219 3939 5225
rect 3881 5185 3893 5219
rect 3927 5216 3939 5219
rect 4154 5216 4160 5228
rect 3927 5188 4160 5216
rect 3927 5185 3939 5188
rect 3881 5179 3939 5185
rect 4154 5176 4160 5188
rect 4212 5176 4218 5228
rect 4614 5176 4620 5228
rect 4672 5176 4678 5228
rect 4724 5225 4752 5256
rect 5460 5256 5701 5284
rect 5460 5228 5488 5256
rect 5689 5253 5701 5256
rect 5735 5253 5747 5287
rect 5689 5247 5747 5253
rect 5902 5244 5908 5296
rect 5960 5244 5966 5296
rect 7561 5287 7619 5293
rect 7561 5253 7573 5287
rect 7607 5284 7619 5287
rect 7760 5284 7788 5315
rect 8294 5312 8300 5324
rect 8352 5352 8358 5364
rect 8662 5352 8668 5364
rect 8352 5324 8668 5352
rect 8352 5312 8358 5324
rect 8662 5312 8668 5324
rect 8720 5312 8726 5364
rect 9214 5312 9220 5364
rect 9272 5352 9278 5364
rect 9272 5324 9674 5352
rect 9272 5312 9278 5324
rect 9646 5284 9674 5324
rect 10318 5312 10324 5364
rect 10376 5352 10382 5364
rect 10965 5355 11023 5361
rect 10965 5352 10977 5355
rect 10376 5324 10977 5352
rect 10376 5312 10382 5324
rect 10965 5321 10977 5324
rect 11011 5321 11023 5355
rect 10965 5315 11023 5321
rect 11698 5312 11704 5364
rect 11756 5352 11762 5364
rect 12529 5355 12587 5361
rect 12529 5352 12541 5355
rect 11756 5324 12541 5352
rect 11756 5312 11762 5324
rect 12529 5321 12541 5324
rect 12575 5321 12587 5355
rect 13722 5352 13728 5364
rect 12529 5315 12587 5321
rect 12636 5324 13728 5352
rect 11146 5284 11152 5296
rect 7607 5256 7788 5284
rect 8036 5256 8616 5284
rect 9646 5256 11152 5284
rect 7607 5253 7619 5256
rect 7561 5247 7619 5253
rect 4709 5219 4767 5225
rect 4709 5185 4721 5219
rect 4755 5216 4767 5219
rect 5169 5219 5227 5225
rect 4755 5188 5120 5216
rect 4755 5185 4767 5188
rect 4709 5179 4767 5185
rect 2869 5151 2927 5157
rect 2869 5117 2881 5151
rect 2915 5148 2927 5151
rect 3973 5151 4031 5157
rect 2915 5120 3556 5148
rect 2915 5117 2927 5120
rect 2869 5111 2927 5117
rect 3528 5089 3556 5120
rect 3973 5117 3985 5151
rect 4019 5148 4031 5151
rect 4341 5151 4399 5157
rect 4341 5148 4353 5151
rect 4019 5120 4353 5148
rect 4019 5117 4031 5120
rect 3973 5111 4031 5117
rect 4341 5117 4353 5120
rect 4387 5117 4399 5151
rect 4632 5148 4660 5176
rect 4985 5151 5043 5157
rect 4985 5148 4997 5151
rect 4632 5120 4997 5148
rect 4341 5111 4399 5117
rect 4985 5117 4997 5120
rect 5031 5117 5043 5151
rect 4985 5111 5043 5117
rect 3513 5083 3571 5089
rect 3513 5049 3525 5083
rect 3559 5049 3571 5083
rect 5092 5080 5120 5188
rect 5169 5185 5181 5219
rect 5215 5185 5227 5219
rect 5169 5179 5227 5185
rect 5184 5148 5212 5179
rect 5442 5176 5448 5228
rect 5500 5176 5506 5228
rect 7190 5176 7196 5228
rect 7248 5176 7254 5228
rect 7466 5176 7472 5228
rect 7524 5216 7530 5228
rect 8036 5216 8064 5256
rect 8588 5225 8616 5256
rect 11146 5244 11152 5256
rect 11204 5244 11210 5296
rect 7524 5188 8064 5216
rect 8573 5219 8631 5225
rect 7524 5176 7530 5188
rect 8573 5185 8585 5219
rect 8619 5185 8631 5219
rect 8573 5179 8631 5185
rect 8757 5219 8815 5225
rect 8757 5185 8769 5219
rect 8803 5216 8815 5219
rect 9122 5216 9128 5228
rect 8803 5188 9128 5216
rect 8803 5185 8815 5188
rect 8757 5179 8815 5185
rect 9122 5176 9128 5188
rect 9180 5176 9186 5228
rect 10134 5176 10140 5228
rect 10192 5216 10198 5228
rect 10229 5219 10287 5225
rect 10229 5216 10241 5219
rect 10192 5188 10241 5216
rect 10192 5176 10198 5188
rect 10229 5185 10241 5188
rect 10275 5185 10287 5219
rect 10229 5179 10287 5185
rect 10410 5176 10416 5228
rect 10468 5176 10474 5228
rect 10502 5176 10508 5228
rect 10560 5216 10566 5228
rect 10597 5219 10655 5225
rect 10597 5216 10609 5219
rect 10560 5188 10609 5216
rect 10560 5176 10566 5188
rect 10597 5185 10609 5188
rect 10643 5185 10655 5219
rect 10597 5179 10655 5185
rect 10686 5176 10692 5228
rect 10744 5176 10750 5228
rect 10778 5176 10784 5228
rect 10836 5176 10842 5228
rect 12636 5216 12664 5324
rect 13722 5312 13728 5324
rect 13780 5312 13786 5364
rect 13814 5312 13820 5364
rect 13872 5352 13878 5364
rect 13872 5324 15424 5352
rect 13872 5312 13878 5324
rect 14090 5284 14096 5296
rect 12728 5256 14096 5284
rect 12728 5225 12756 5256
rect 14090 5244 14096 5256
rect 14148 5244 14154 5296
rect 12452 5188 12664 5216
rect 12713 5219 12771 5225
rect 5902 5148 5908 5160
rect 5184 5120 5908 5148
rect 5902 5108 5908 5120
rect 5960 5108 5966 5160
rect 7374 5108 7380 5160
rect 7432 5108 7438 5160
rect 7650 5108 7656 5160
rect 7708 5148 7714 5160
rect 8205 5151 8263 5157
rect 8205 5148 8217 5151
rect 7708 5120 8217 5148
rect 7708 5108 7714 5120
rect 8205 5117 8217 5120
rect 8251 5117 8263 5151
rect 8205 5111 8263 5117
rect 8389 5151 8447 5157
rect 8389 5117 8401 5151
rect 8435 5148 8447 5151
rect 9214 5148 9220 5160
rect 8435 5120 9220 5148
rect 8435 5117 8447 5120
rect 8389 5111 8447 5117
rect 9214 5108 9220 5120
rect 9272 5108 9278 5160
rect 9490 5108 9496 5160
rect 9548 5148 9554 5160
rect 12452 5148 12480 5188
rect 12713 5185 12725 5219
rect 12759 5185 12771 5219
rect 12713 5179 12771 5185
rect 12802 5176 12808 5228
rect 12860 5176 12866 5228
rect 13081 5219 13139 5225
rect 13081 5185 13093 5219
rect 13127 5185 13139 5219
rect 13081 5179 13139 5185
rect 9548 5120 12480 5148
rect 9548 5108 9554 5120
rect 12526 5108 12532 5160
rect 12584 5148 12590 5160
rect 13096 5148 13124 5179
rect 14274 5176 14280 5228
rect 14332 5176 14338 5228
rect 14366 5176 14372 5228
rect 14424 5176 14430 5228
rect 14550 5176 14556 5228
rect 14608 5216 14614 5228
rect 15286 5225 15292 5228
rect 14645 5219 14703 5225
rect 14645 5216 14657 5219
rect 14608 5188 14657 5216
rect 14608 5176 14614 5188
rect 14645 5185 14657 5188
rect 14691 5185 14703 5219
rect 15277 5219 15292 5225
rect 15277 5216 15289 5219
rect 14645 5179 14703 5185
rect 14752 5188 15289 5216
rect 12584 5120 13124 5148
rect 12584 5108 12590 5120
rect 13722 5108 13728 5160
rect 13780 5148 13786 5160
rect 14752 5148 14780 5188
rect 15277 5185 15289 5188
rect 15277 5179 15292 5185
rect 15286 5176 15292 5179
rect 15344 5176 15350 5228
rect 15396 5216 15424 5324
rect 16298 5312 16304 5364
rect 16356 5352 16362 5364
rect 16393 5355 16451 5361
rect 16393 5352 16405 5355
rect 16356 5324 16405 5352
rect 16356 5312 16362 5324
rect 16393 5321 16405 5324
rect 16439 5321 16451 5355
rect 16393 5315 16451 5321
rect 15930 5244 15936 5296
rect 15988 5284 15994 5296
rect 15988 5256 16712 5284
rect 15988 5244 15994 5256
rect 15473 5219 15531 5225
rect 15473 5216 15485 5219
rect 15396 5188 15485 5216
rect 15473 5185 15485 5188
rect 15519 5185 15531 5219
rect 15473 5179 15531 5185
rect 16022 5176 16028 5228
rect 16080 5176 16086 5228
rect 16684 5225 16712 5256
rect 16669 5219 16727 5225
rect 16669 5185 16681 5219
rect 16715 5185 16727 5219
rect 16669 5179 16727 5185
rect 16853 5219 16911 5225
rect 16853 5185 16865 5219
rect 16899 5185 16911 5219
rect 16853 5179 16911 5185
rect 13780 5120 14780 5148
rect 15381 5151 15439 5157
rect 13780 5108 13786 5120
rect 15381 5117 15393 5151
rect 15427 5148 15439 5151
rect 16117 5151 16175 5157
rect 16117 5148 16129 5151
rect 15427 5120 16129 5148
rect 15427 5117 15439 5120
rect 15381 5111 15439 5117
rect 16117 5117 16129 5120
rect 16163 5148 16175 5151
rect 16868 5148 16896 5179
rect 16163 5120 16896 5148
rect 16163 5117 16175 5120
rect 16117 5111 16175 5117
rect 5537 5083 5595 5089
rect 5537 5080 5549 5083
rect 5092 5052 5549 5080
rect 3513 5043 3571 5049
rect 5537 5049 5549 5052
rect 5583 5049 5595 5083
rect 5537 5043 5595 5049
rect 7190 5040 7196 5092
rect 7248 5040 7254 5092
rect 10045 5083 10103 5089
rect 10045 5080 10057 5083
rect 8588 5052 10057 5080
rect 5721 5015 5779 5021
rect 5721 4981 5733 5015
rect 5767 5012 5779 5015
rect 5810 5012 5816 5024
rect 5767 4984 5816 5012
rect 5767 4981 5779 4984
rect 5721 4975 5779 4981
rect 5810 4972 5816 4984
rect 5868 5012 5874 5024
rect 6638 5012 6644 5024
rect 5868 4984 6644 5012
rect 5868 4972 5874 4984
rect 6638 4972 6644 4984
rect 6696 5012 6702 5024
rect 8588 5012 8616 5052
rect 10045 5049 10057 5052
rect 10091 5049 10103 5083
rect 10045 5043 10103 5049
rect 10962 5040 10968 5092
rect 11020 5080 11026 5092
rect 14093 5083 14151 5089
rect 14093 5080 14105 5083
rect 11020 5052 14105 5080
rect 11020 5040 11026 5052
rect 14093 5049 14105 5052
rect 14139 5049 14151 5083
rect 14093 5043 14151 5049
rect 6696 4984 8616 5012
rect 6696 4972 6702 4984
rect 8662 4972 8668 5024
rect 8720 5012 8726 5024
rect 9306 5012 9312 5024
rect 8720 4984 9312 5012
rect 8720 4972 8726 4984
rect 9306 4972 9312 4984
rect 9364 4972 9370 5024
rect 10226 4972 10232 5024
rect 10284 4972 10290 5024
rect 12894 4972 12900 5024
rect 12952 5012 12958 5024
rect 12989 5015 13047 5021
rect 12989 5012 13001 5015
rect 12952 4984 13001 5012
rect 12952 4972 12958 4984
rect 12989 4981 13001 4984
rect 13035 5012 13047 5015
rect 14550 5012 14556 5024
rect 13035 4984 14556 5012
rect 13035 4981 13047 4984
rect 12989 4975 13047 4981
rect 14550 4972 14556 4984
rect 14608 4972 14614 5024
rect 15930 4972 15936 5024
rect 15988 5012 15994 5024
rect 16025 5015 16083 5021
rect 16025 5012 16037 5015
rect 15988 4984 16037 5012
rect 15988 4972 15994 4984
rect 16025 4981 16037 4984
rect 16071 4981 16083 5015
rect 16025 4975 16083 4981
rect 16669 5015 16727 5021
rect 16669 4981 16681 5015
rect 16715 5012 16727 5015
rect 16758 5012 16764 5024
rect 16715 4984 16764 5012
rect 16715 4981 16727 4984
rect 16669 4975 16727 4981
rect 16758 4972 16764 4984
rect 16816 4972 16822 5024
rect 1104 4922 17848 4944
rect 1104 4870 1918 4922
rect 1970 4870 1982 4922
rect 2034 4870 2046 4922
rect 2098 4870 2110 4922
rect 2162 4870 2174 4922
rect 2226 4870 2238 4922
rect 2290 4870 7918 4922
rect 7970 4870 7982 4922
rect 8034 4870 8046 4922
rect 8098 4870 8110 4922
rect 8162 4870 8174 4922
rect 8226 4870 8238 4922
rect 8290 4870 13918 4922
rect 13970 4870 13982 4922
rect 14034 4870 14046 4922
rect 14098 4870 14110 4922
rect 14162 4870 14174 4922
rect 14226 4870 14238 4922
rect 14290 4870 17848 4922
rect 1104 4848 17848 4870
rect 2314 4768 2320 4820
rect 2372 4768 2378 4820
rect 5442 4768 5448 4820
rect 5500 4808 5506 4820
rect 10042 4808 10048 4820
rect 5500 4780 10048 4808
rect 5500 4768 5506 4780
rect 10042 4768 10048 4780
rect 10100 4768 10106 4820
rect 10686 4768 10692 4820
rect 10744 4808 10750 4820
rect 10873 4811 10931 4817
rect 10873 4808 10885 4811
rect 10744 4780 10885 4808
rect 10744 4768 10750 4780
rect 10873 4777 10885 4780
rect 10919 4777 10931 4811
rect 10873 4771 10931 4777
rect 11241 4811 11299 4817
rect 11241 4777 11253 4811
rect 11287 4808 11299 4811
rect 12250 4808 12256 4820
rect 11287 4780 12256 4808
rect 11287 4777 11299 4780
rect 11241 4771 11299 4777
rect 12250 4768 12256 4780
rect 12308 4768 12314 4820
rect 16574 4768 16580 4820
rect 16632 4808 16638 4820
rect 16761 4811 16819 4817
rect 16761 4808 16773 4811
rect 16632 4780 16773 4808
rect 16632 4768 16638 4780
rect 16761 4777 16773 4780
rect 16807 4777 16819 4811
rect 16761 4771 16819 4777
rect 8386 4700 8392 4752
rect 8444 4740 8450 4752
rect 9122 4740 9128 4752
rect 8444 4712 9128 4740
rect 8444 4700 8450 4712
rect 9122 4700 9128 4712
rect 9180 4700 9186 4752
rect 9677 4743 9735 4749
rect 9677 4709 9689 4743
rect 9723 4740 9735 4743
rect 10502 4740 10508 4752
rect 9723 4712 10508 4740
rect 9723 4709 9735 4712
rect 9677 4703 9735 4709
rect 7558 4632 7564 4684
rect 7616 4672 7622 4684
rect 7616 4644 9168 4672
rect 7616 4632 7622 4644
rect 1578 4564 1584 4616
rect 1636 4564 1642 4616
rect 2406 4564 2412 4616
rect 2464 4564 2470 4616
rect 6181 4607 6239 4613
rect 6181 4573 6193 4607
rect 6227 4573 6239 4607
rect 6181 4567 6239 4573
rect 6196 4536 6224 4567
rect 6362 4564 6368 4616
rect 6420 4564 6426 4616
rect 8570 4564 8576 4616
rect 8628 4604 8634 4616
rect 9140 4613 9168 4644
rect 9306 4632 9312 4684
rect 9364 4632 9370 4684
rect 10152 4681 10180 4712
rect 10502 4700 10508 4712
rect 10560 4700 10566 4752
rect 10137 4675 10195 4681
rect 10137 4641 10149 4675
rect 10183 4641 10195 4675
rect 10137 4635 10195 4641
rect 10597 4675 10655 4681
rect 10597 4641 10609 4675
rect 10643 4672 10655 4675
rect 10704 4672 10732 4768
rect 16666 4700 16672 4752
rect 16724 4700 16730 4752
rect 16853 4743 16911 4749
rect 16853 4709 16865 4743
rect 16899 4709 16911 4743
rect 16853 4703 16911 4709
rect 10643 4644 10732 4672
rect 10781 4675 10839 4681
rect 10643 4641 10655 4644
rect 10597 4635 10655 4641
rect 10781 4641 10793 4675
rect 10827 4672 10839 4675
rect 10870 4672 10876 4684
rect 10827 4644 10876 4672
rect 10827 4641 10839 4644
rect 10781 4635 10839 4641
rect 10870 4632 10876 4644
rect 10928 4632 10934 4684
rect 11146 4632 11152 4684
rect 11204 4672 11210 4684
rect 11606 4672 11612 4684
rect 11204 4644 11612 4672
rect 11204 4632 11210 4644
rect 11606 4632 11612 4644
rect 11664 4632 11670 4684
rect 15562 4632 15568 4684
rect 15620 4672 15626 4684
rect 16022 4672 16028 4684
rect 15620 4644 16028 4672
rect 15620 4632 15626 4644
rect 16022 4632 16028 4644
rect 16080 4672 16086 4684
rect 16209 4675 16267 4681
rect 16209 4672 16221 4675
rect 16080 4644 16221 4672
rect 16080 4632 16086 4644
rect 16209 4641 16221 4644
rect 16255 4672 16267 4675
rect 16868 4672 16896 4703
rect 16255 4644 16896 4672
rect 16255 4641 16267 4644
rect 16209 4635 16267 4641
rect 8941 4607 8999 4613
rect 8941 4604 8953 4607
rect 8628 4576 8953 4604
rect 8628 4564 8634 4576
rect 8941 4573 8953 4576
rect 8987 4573 8999 4607
rect 8941 4567 8999 4573
rect 9125 4607 9183 4613
rect 9125 4573 9137 4607
rect 9171 4573 9183 4607
rect 9125 4567 9183 4573
rect 7190 4536 7196 4548
rect 6196 4508 7196 4536
rect 7190 4496 7196 4508
rect 7248 4496 7254 4548
rect 842 4428 848 4480
rect 900 4468 906 4480
rect 1397 4471 1455 4477
rect 1397 4468 1409 4471
rect 900 4440 1409 4468
rect 900 4428 906 4440
rect 1397 4437 1409 4440
rect 1443 4437 1455 4471
rect 1397 4431 1455 4437
rect 6178 4428 6184 4480
rect 6236 4428 6242 4480
rect 7098 4428 7104 4480
rect 7156 4468 7162 4480
rect 7650 4468 7656 4480
rect 7156 4440 7656 4468
rect 7156 4428 7162 4440
rect 7650 4428 7656 4440
rect 7708 4428 7714 4480
rect 9140 4468 9168 4567
rect 9214 4564 9220 4616
rect 9272 4564 9278 4616
rect 9490 4564 9496 4616
rect 9548 4564 9554 4616
rect 10505 4607 10563 4613
rect 10505 4573 10517 4607
rect 10551 4604 10563 4607
rect 10686 4604 10692 4616
rect 10551 4576 10692 4604
rect 10551 4573 10563 4576
rect 10505 4567 10563 4573
rect 10686 4564 10692 4576
rect 10744 4564 10750 4616
rect 11241 4607 11299 4613
rect 11241 4573 11253 4607
rect 11287 4604 11299 4607
rect 11422 4604 11428 4616
rect 11287 4576 11428 4604
rect 11287 4573 11299 4576
rect 11241 4567 11299 4573
rect 11422 4564 11428 4576
rect 11480 4564 11486 4616
rect 16301 4607 16359 4613
rect 16301 4573 16313 4607
rect 16347 4604 16359 4607
rect 16758 4604 16764 4616
rect 16347 4576 16764 4604
rect 16347 4573 16359 4576
rect 16301 4567 16359 4573
rect 16758 4564 16764 4576
rect 16816 4604 16822 4616
rect 17221 4607 17279 4613
rect 17221 4604 17233 4607
rect 16816 4576 17233 4604
rect 16816 4564 16822 4576
rect 17221 4573 17233 4576
rect 17267 4573 17279 4607
rect 17221 4567 17279 4573
rect 9232 4536 9260 4564
rect 13354 4536 13360 4548
rect 9232 4508 13360 4536
rect 13354 4496 13360 4508
rect 13412 4496 13418 4548
rect 13814 4468 13820 4480
rect 9140 4440 13820 4468
rect 13814 4428 13820 4440
rect 13872 4428 13878 4480
rect 1104 4378 17848 4400
rect 1104 4326 2658 4378
rect 2710 4326 2722 4378
rect 2774 4326 2786 4378
rect 2838 4326 2850 4378
rect 2902 4326 2914 4378
rect 2966 4326 2978 4378
rect 3030 4326 8658 4378
rect 8710 4326 8722 4378
rect 8774 4326 8786 4378
rect 8838 4326 8850 4378
rect 8902 4326 8914 4378
rect 8966 4326 8978 4378
rect 9030 4326 14658 4378
rect 14710 4326 14722 4378
rect 14774 4326 14786 4378
rect 14838 4326 14850 4378
rect 14902 4326 14914 4378
rect 14966 4326 14978 4378
rect 15030 4326 17848 4378
rect 1104 4304 17848 4326
rect 4154 4224 4160 4276
rect 4212 4264 4218 4276
rect 4341 4267 4399 4273
rect 4341 4264 4353 4267
rect 4212 4236 4353 4264
rect 4212 4224 4218 4236
rect 4341 4233 4353 4236
rect 4387 4233 4399 4267
rect 4341 4227 4399 4233
rect 8570 4224 8576 4276
rect 8628 4264 8634 4276
rect 8665 4267 8723 4273
rect 8665 4264 8677 4267
rect 8628 4236 8677 4264
rect 8628 4224 8634 4236
rect 8665 4233 8677 4236
rect 8711 4233 8723 4267
rect 8665 4227 8723 4233
rect 10870 4224 10876 4276
rect 10928 4264 10934 4276
rect 11057 4267 11115 4273
rect 11057 4264 11069 4267
rect 10928 4236 11069 4264
rect 10928 4224 10934 4236
rect 11057 4233 11069 4236
rect 11103 4264 11115 4267
rect 11238 4264 11244 4276
rect 11103 4236 11244 4264
rect 11103 4233 11115 4236
rect 11057 4227 11115 4233
rect 11238 4224 11244 4236
rect 11296 4264 11302 4276
rect 11974 4264 11980 4276
rect 11296 4236 11980 4264
rect 11296 4224 11302 4236
rect 11974 4224 11980 4236
rect 12032 4224 12038 4276
rect 12342 4224 12348 4276
rect 12400 4224 12406 4276
rect 12434 4224 12440 4276
rect 12492 4264 12498 4276
rect 12713 4267 12771 4273
rect 12713 4264 12725 4267
rect 12492 4236 12725 4264
rect 12492 4224 12498 4236
rect 12713 4233 12725 4236
rect 12759 4233 12771 4267
rect 12713 4227 12771 4233
rect 13446 4224 13452 4276
rect 13504 4224 13510 4276
rect 14826 4224 14832 4276
rect 14884 4224 14890 4276
rect 3329 4199 3387 4205
rect 3329 4196 3341 4199
rect 2438 4168 3341 4196
rect 3329 4165 3341 4168
rect 3375 4165 3387 4199
rect 3329 4159 3387 4165
rect 5905 4199 5963 4205
rect 5905 4165 5917 4199
rect 5951 4196 5963 4199
rect 7101 4199 7159 4205
rect 7101 4196 7113 4199
rect 5951 4168 7113 4196
rect 5951 4165 5963 4168
rect 5905 4159 5963 4165
rect 7101 4165 7113 4168
rect 7147 4165 7159 4199
rect 7101 4159 7159 4165
rect 11422 4156 11428 4208
rect 11480 4196 11486 4208
rect 12360 4196 12388 4224
rect 11480 4168 12756 4196
rect 11480 4156 11486 4168
rect 3142 4088 3148 4140
rect 3200 4088 3206 4140
rect 3421 4131 3479 4137
rect 3421 4097 3433 4131
rect 3467 4128 3479 4131
rect 3510 4128 3516 4140
rect 3467 4100 3516 4128
rect 3467 4097 3479 4100
rect 3421 4091 3479 4097
rect 3510 4088 3516 4100
rect 3568 4088 3574 4140
rect 4065 4131 4123 4137
rect 4065 4097 4077 4131
rect 4111 4128 4123 4131
rect 4111 4100 4844 4128
rect 4111 4097 4123 4100
rect 4065 4091 4123 4097
rect 1397 4063 1455 4069
rect 1397 4029 1409 4063
rect 1443 4060 1455 4063
rect 1486 4060 1492 4072
rect 1443 4032 1492 4060
rect 1443 4029 1455 4032
rect 1397 4023 1455 4029
rect 1486 4020 1492 4032
rect 1544 4020 1550 4072
rect 4816 4069 4844 4100
rect 6086 4088 6092 4140
rect 6144 4088 6150 4140
rect 6178 4088 6184 4140
rect 6236 4088 6242 4140
rect 6733 4131 6791 4137
rect 6733 4097 6745 4131
rect 6779 4128 6791 4131
rect 6914 4128 6920 4140
rect 6779 4100 6920 4128
rect 6779 4097 6791 4100
rect 6733 4091 6791 4097
rect 6914 4088 6920 4100
rect 6972 4088 6978 4140
rect 7009 4131 7067 4137
rect 7009 4097 7021 4131
rect 7055 4097 7067 4131
rect 7009 4091 7067 4097
rect 2869 4063 2927 4069
rect 2869 4029 2881 4063
rect 2915 4060 2927 4063
rect 4157 4063 4215 4069
rect 2915 4032 3740 4060
rect 2915 4029 2927 4032
rect 2869 4023 2927 4029
rect 3712 4001 3740 4032
rect 4157 4029 4169 4063
rect 4203 4029 4215 4063
rect 4157 4023 4215 4029
rect 4801 4063 4859 4069
rect 4801 4029 4813 4063
rect 4847 4060 4859 4063
rect 4847 4032 6040 4060
rect 4847 4029 4859 4032
rect 4801 4023 4859 4029
rect 3697 3995 3755 4001
rect 3697 3961 3709 3995
rect 3743 3961 3755 3995
rect 4172 3992 4200 4023
rect 4522 3992 4528 4004
rect 4172 3964 4528 3992
rect 3697 3955 3755 3961
rect 4522 3952 4528 3964
rect 4580 3952 4586 4004
rect 5902 3952 5908 4004
rect 5960 3952 5966 4004
rect 6012 3992 6040 4032
rect 6362 4020 6368 4072
rect 6420 4060 6426 4072
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6420 4032 6837 4060
rect 6420 4020 6426 4032
rect 6825 4029 6837 4032
rect 6871 4060 6883 4063
rect 7024 4060 7052 4091
rect 7190 4088 7196 4140
rect 7248 4088 7254 4140
rect 7466 4088 7472 4140
rect 7524 4128 7530 4140
rect 8297 4131 8355 4137
rect 8297 4128 8309 4131
rect 7524 4100 8309 4128
rect 7524 4088 7530 4100
rect 8297 4097 8309 4100
rect 8343 4097 8355 4131
rect 8297 4091 8355 4097
rect 6871 4032 7052 4060
rect 8312 4060 8340 4091
rect 8386 4088 8392 4140
rect 8444 4088 8450 4140
rect 8481 4131 8539 4137
rect 8481 4097 8493 4131
rect 8527 4128 8539 4131
rect 9490 4128 9496 4140
rect 8527 4100 9496 4128
rect 8527 4097 8539 4100
rect 8481 4091 8539 4097
rect 9490 4088 9496 4100
rect 9548 4088 9554 4140
rect 10796 4100 12204 4128
rect 8662 4060 8668 4072
rect 8312 4032 8668 4060
rect 6871 4029 6883 4032
rect 6825 4023 6883 4029
rect 6546 3992 6552 4004
rect 6012 3964 6552 3992
rect 6546 3952 6552 3964
rect 6604 3952 6610 4004
rect 6362 3884 6368 3936
rect 6420 3924 6426 3936
rect 6457 3927 6515 3933
rect 6457 3924 6469 3927
rect 6420 3896 6469 3924
rect 6420 3884 6426 3896
rect 6457 3893 6469 3896
rect 6503 3893 6515 3927
rect 7024 3924 7052 4032
rect 8662 4020 8668 4032
rect 8720 4020 8726 4072
rect 10796 4004 10824 4100
rect 12069 4063 12127 4069
rect 12069 4060 12081 4063
rect 10888 4032 12081 4060
rect 7650 3952 7656 4004
rect 7708 3992 7714 4004
rect 10689 3995 10747 4001
rect 10689 3992 10701 3995
rect 7708 3964 10701 3992
rect 7708 3952 7714 3964
rect 10689 3961 10701 3964
rect 10735 3992 10747 3995
rect 10778 3992 10784 4004
rect 10735 3964 10784 3992
rect 10735 3961 10747 3964
rect 10689 3955 10747 3961
rect 10778 3952 10784 3964
rect 10836 3952 10842 4004
rect 10888 3924 10916 4032
rect 12069 4029 12081 4032
rect 12115 4029 12127 4063
rect 12176 4060 12204 4100
rect 12250 4088 12256 4140
rect 12308 4088 12314 4140
rect 12434 4137 12440 4140
rect 12391 4131 12440 4137
rect 12391 4129 12403 4131
rect 12348 4101 12403 4129
rect 12391 4097 12403 4101
rect 12437 4097 12440 4131
rect 12391 4091 12440 4097
rect 12434 4088 12440 4091
rect 12492 4088 12498 4140
rect 12621 4131 12679 4137
rect 12621 4097 12633 4131
rect 12667 4097 12679 4131
rect 12728 4128 12756 4168
rect 12802 4156 12808 4208
rect 12860 4196 12866 4208
rect 13357 4199 13415 4205
rect 12860 4168 13124 4196
rect 12860 4156 12866 4168
rect 12989 4131 13047 4137
rect 12989 4128 13001 4131
rect 12728 4100 13001 4128
rect 12621 4091 12679 4097
rect 12989 4097 13001 4100
rect 13035 4097 13047 4131
rect 13096 4128 13124 4168
rect 13357 4165 13369 4199
rect 13403 4196 13415 4199
rect 13464 4196 13492 4224
rect 14458 4196 14464 4208
rect 13403 4168 13492 4196
rect 13832 4168 14464 4196
rect 13403 4165 13415 4168
rect 13357 4159 13415 4165
rect 13265 4131 13323 4137
rect 13265 4128 13277 4131
rect 13096 4100 13277 4128
rect 12989 4091 13047 4097
rect 13265 4097 13277 4100
rect 13311 4097 13323 4131
rect 13265 4091 13323 4097
rect 12636 4060 12664 4091
rect 13538 4088 13544 4140
rect 13596 4128 13602 4140
rect 13832 4137 13860 4168
rect 14458 4156 14464 4168
rect 14516 4196 14522 4208
rect 15838 4196 15844 4208
rect 14516 4168 15844 4196
rect 14516 4156 14522 4168
rect 15838 4156 15844 4168
rect 15896 4156 15902 4208
rect 13725 4131 13783 4137
rect 13725 4128 13737 4131
rect 13596 4100 13737 4128
rect 13596 4088 13602 4100
rect 13725 4097 13737 4100
rect 13771 4097 13783 4131
rect 13725 4091 13783 4097
rect 13817 4131 13875 4137
rect 13817 4097 13829 4131
rect 13863 4097 13875 4131
rect 13817 4091 13875 4097
rect 12897 4063 12955 4069
rect 12897 4060 12909 4063
rect 12176 4032 12909 4060
rect 12069 4023 12127 4029
rect 12897 4029 12909 4032
rect 12943 4029 12955 4063
rect 12897 4023 12955 4029
rect 13630 4020 13636 4072
rect 13688 4020 13694 4072
rect 12434 3952 12440 4004
rect 12492 3992 12498 4004
rect 13832 3992 13860 4091
rect 14366 4088 14372 4140
rect 14424 4128 14430 4140
rect 14770 4131 14828 4137
rect 14770 4128 14782 4131
rect 14424 4100 14782 4128
rect 14424 4088 14430 4100
rect 14770 4097 14782 4100
rect 14816 4097 14828 4131
rect 15565 4131 15623 4137
rect 15565 4128 15577 4131
rect 14770 4091 14828 4097
rect 14936 4100 15577 4128
rect 14936 4060 14964 4100
rect 15565 4097 15577 4100
rect 15611 4097 15623 4131
rect 15565 4091 15623 4097
rect 15657 4131 15715 4137
rect 15657 4097 15669 4131
rect 15703 4128 15715 4131
rect 15746 4128 15752 4140
rect 15703 4100 15752 4128
rect 15703 4097 15715 4100
rect 15657 4091 15715 4097
rect 15746 4088 15752 4100
rect 15804 4088 15810 4140
rect 12492 3964 13860 3992
rect 13924 4032 14964 4060
rect 12492 3952 12498 3964
rect 7024 3896 10916 3924
rect 11057 3927 11115 3933
rect 6457 3887 6515 3893
rect 11057 3893 11069 3927
rect 11103 3924 11115 3927
rect 11146 3924 11152 3936
rect 11103 3896 11152 3924
rect 11103 3893 11115 3896
rect 11057 3887 11115 3893
rect 11146 3884 11152 3896
rect 11204 3884 11210 3936
rect 11238 3884 11244 3936
rect 11296 3884 11302 3936
rect 12529 3927 12587 3933
rect 12529 3893 12541 3927
rect 12575 3924 12587 3927
rect 12894 3924 12900 3936
rect 12575 3896 12900 3924
rect 12575 3893 12587 3896
rect 12529 3887 12587 3893
rect 12894 3884 12900 3896
rect 12952 3884 12958 3936
rect 13722 3884 13728 3936
rect 13780 3924 13786 3936
rect 13924 3924 13952 4032
rect 15286 4020 15292 4072
rect 15344 4020 15350 4072
rect 15378 4020 15384 4072
rect 15436 4020 15442 4072
rect 14645 3995 14703 4001
rect 14645 3961 14657 3995
rect 14691 3992 14703 3995
rect 15102 3992 15108 4004
rect 14691 3964 15108 3992
rect 14691 3961 14703 3964
rect 14645 3955 14703 3961
rect 15102 3952 15108 3964
rect 15160 3952 15166 4004
rect 13780 3896 13952 3924
rect 13780 3884 13786 3896
rect 14550 3884 14556 3936
rect 14608 3924 14614 3936
rect 15197 3927 15255 3933
rect 15197 3924 15209 3927
rect 14608 3896 15209 3924
rect 14608 3884 14614 3896
rect 15197 3893 15209 3896
rect 15243 3893 15255 3927
rect 15197 3887 15255 3893
rect 15470 3884 15476 3936
rect 15528 3884 15534 3936
rect 1104 3834 17848 3856
rect 1104 3782 1918 3834
rect 1970 3782 1982 3834
rect 2034 3782 2046 3834
rect 2098 3782 2110 3834
rect 2162 3782 2174 3834
rect 2226 3782 2238 3834
rect 2290 3782 7918 3834
rect 7970 3782 7982 3834
rect 8034 3782 8046 3834
rect 8098 3782 8110 3834
rect 8162 3782 8174 3834
rect 8226 3782 8238 3834
rect 8290 3782 13918 3834
rect 13970 3782 13982 3834
rect 14034 3782 14046 3834
rect 14098 3782 14110 3834
rect 14162 3782 14174 3834
rect 14226 3782 14238 3834
rect 14290 3782 17848 3834
rect 1104 3760 17848 3782
rect 4522 3680 4528 3732
rect 4580 3720 4586 3732
rect 5905 3723 5963 3729
rect 5905 3720 5917 3723
rect 4580 3692 5917 3720
rect 4580 3680 4586 3692
rect 5905 3689 5917 3692
rect 5951 3689 5963 3723
rect 5905 3683 5963 3689
rect 8294 3680 8300 3732
rect 8352 3680 8358 3732
rect 8481 3723 8539 3729
rect 8481 3689 8493 3723
rect 8527 3689 8539 3723
rect 8481 3683 8539 3689
rect 3436 3624 6500 3652
rect 3436 3593 3464 3624
rect 3421 3587 3479 3593
rect 3421 3553 3433 3587
rect 3467 3553 3479 3587
rect 3421 3547 3479 3553
rect 6362 3544 6368 3596
rect 6420 3544 6426 3596
rect 6472 3584 6500 3624
rect 6546 3612 6552 3664
rect 6604 3652 6610 3664
rect 7837 3655 7895 3661
rect 7837 3652 7849 3655
rect 6604 3624 7849 3652
rect 6604 3612 6610 3624
rect 7837 3621 7849 3624
rect 7883 3621 7895 3655
rect 8386 3652 8392 3664
rect 7837 3615 7895 3621
rect 7944 3624 8392 3652
rect 7944 3584 7972 3624
rect 8386 3612 8392 3624
rect 8444 3612 8450 3664
rect 8496 3652 8524 3683
rect 10686 3680 10692 3732
rect 10744 3680 10750 3732
rect 12250 3680 12256 3732
rect 12308 3720 12314 3732
rect 12989 3723 13047 3729
rect 12989 3720 13001 3723
rect 12308 3692 13001 3720
rect 12308 3680 12314 3692
rect 12989 3689 13001 3692
rect 13035 3689 13047 3723
rect 12989 3683 13047 3689
rect 13170 3680 13176 3732
rect 13228 3720 13234 3732
rect 13357 3723 13415 3729
rect 13357 3720 13369 3723
rect 13228 3692 13369 3720
rect 13228 3680 13234 3692
rect 13357 3689 13369 3692
rect 13403 3720 13415 3723
rect 13722 3720 13728 3732
rect 13403 3692 13728 3720
rect 13403 3689 13415 3692
rect 13357 3683 13415 3689
rect 13722 3680 13728 3692
rect 13780 3680 13786 3732
rect 13817 3723 13875 3729
rect 13817 3689 13829 3723
rect 13863 3720 13875 3723
rect 14366 3720 14372 3732
rect 13863 3692 14372 3720
rect 13863 3689 13875 3692
rect 13817 3683 13875 3689
rect 14366 3680 14372 3692
rect 14424 3680 14430 3732
rect 14550 3680 14556 3732
rect 14608 3720 14614 3732
rect 14608 3692 14780 3720
rect 14608 3680 14614 3692
rect 12710 3652 12716 3664
rect 8496 3624 12716 3652
rect 12710 3612 12716 3624
rect 12768 3612 12774 3664
rect 12894 3612 12900 3664
rect 12952 3652 12958 3664
rect 13538 3652 13544 3664
rect 12952 3624 13544 3652
rect 12952 3612 12958 3624
rect 13538 3612 13544 3624
rect 13596 3612 13602 3664
rect 14752 3652 14780 3692
rect 14826 3680 14832 3732
rect 14884 3680 14890 3732
rect 15562 3680 15568 3732
rect 15620 3680 15626 3732
rect 15013 3655 15071 3661
rect 15013 3652 15025 3655
rect 14752 3624 15025 3652
rect 15013 3621 15025 3624
rect 15059 3652 15071 3655
rect 16025 3655 16083 3661
rect 16025 3652 16037 3655
rect 15059 3624 16037 3652
rect 15059 3621 15071 3624
rect 15013 3615 15071 3621
rect 16025 3621 16037 3624
rect 16071 3621 16083 3655
rect 16025 3615 16083 3621
rect 8294 3584 8300 3596
rect 6472 3556 7972 3584
rect 8128 3556 8300 3584
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3516 1639 3519
rect 1627 3488 2774 3516
rect 1627 3485 1639 3488
rect 1581 3479 1639 3485
rect 2746 3448 2774 3488
rect 3234 3476 3240 3528
rect 3292 3476 3298 3528
rect 6086 3476 6092 3528
rect 6144 3516 6150 3528
rect 7484 3525 7512 3556
rect 6273 3519 6331 3525
rect 6273 3516 6285 3519
rect 6144 3488 6285 3516
rect 6144 3476 6150 3488
rect 6273 3485 6285 3488
rect 6319 3485 6331 3519
rect 6273 3479 6331 3485
rect 7469 3519 7527 3525
rect 7469 3485 7481 3519
rect 7515 3485 7527 3519
rect 7469 3479 7527 3485
rect 4246 3448 4252 3460
rect 2746 3420 4252 3448
rect 4246 3408 4252 3420
rect 4304 3408 4310 3460
rect 842 3340 848 3392
rect 900 3380 906 3392
rect 1397 3383 1455 3389
rect 1397 3380 1409 3383
rect 900 3352 1409 3380
rect 900 3340 906 3352
rect 1397 3349 1409 3352
rect 1443 3349 1455 3383
rect 1397 3343 1455 3349
rect 3053 3383 3111 3389
rect 3053 3349 3065 3383
rect 3099 3380 3111 3383
rect 3878 3380 3884 3392
rect 3099 3352 3884 3380
rect 3099 3349 3111 3352
rect 3053 3343 3111 3349
rect 3878 3340 3884 3352
rect 3936 3340 3942 3392
rect 6288 3380 6316 3479
rect 7650 3476 7656 3528
rect 7708 3476 7714 3528
rect 8128 3525 8156 3556
rect 8294 3544 8300 3556
rect 8352 3544 8358 3596
rect 8478 3544 8484 3596
rect 8536 3584 8542 3596
rect 9217 3587 9275 3593
rect 9217 3584 9229 3587
rect 8536 3556 9229 3584
rect 8536 3544 8542 3556
rect 9217 3553 9229 3556
rect 9263 3553 9275 3587
rect 9217 3547 9275 3553
rect 9309 3587 9367 3593
rect 9309 3553 9321 3587
rect 9355 3584 9367 3587
rect 9766 3584 9772 3596
rect 9355 3556 9772 3584
rect 9355 3553 9367 3556
rect 9309 3547 9367 3553
rect 9766 3544 9772 3556
rect 9824 3544 9830 3596
rect 11149 3587 11207 3593
rect 11149 3553 11161 3587
rect 11195 3584 11207 3587
rect 11698 3584 11704 3596
rect 11195 3556 11704 3584
rect 11195 3553 11207 3556
rect 11149 3547 11207 3553
rect 11698 3544 11704 3556
rect 11756 3544 11762 3596
rect 12158 3544 12164 3596
rect 12216 3584 12222 3596
rect 12253 3587 12311 3593
rect 12253 3584 12265 3587
rect 12216 3556 12265 3584
rect 12216 3544 12222 3556
rect 12253 3553 12265 3556
rect 12299 3584 12311 3587
rect 13909 3587 13967 3593
rect 13909 3584 13921 3587
rect 12299 3556 13921 3584
rect 12299 3553 12311 3556
rect 12253 3547 12311 3553
rect 8112 3519 8170 3525
rect 8112 3485 8124 3519
rect 8158 3485 8170 3519
rect 8112 3479 8170 3485
rect 8205 3519 8263 3525
rect 8205 3485 8217 3519
rect 8251 3516 8263 3519
rect 8496 3516 8524 3544
rect 8251 3488 8524 3516
rect 9125 3519 9183 3525
rect 8251 3485 8263 3488
rect 8205 3479 8263 3485
rect 9125 3485 9137 3519
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 7098 3408 7104 3460
rect 7156 3448 7162 3460
rect 7561 3451 7619 3457
rect 7561 3448 7573 3451
rect 7156 3420 7573 3448
rect 7156 3408 7162 3420
rect 7561 3417 7573 3420
rect 7607 3448 7619 3451
rect 8449 3451 8507 3457
rect 8449 3448 8461 3451
rect 7607 3420 8461 3448
rect 7607 3417 7619 3420
rect 7561 3411 7619 3417
rect 8449 3417 8461 3420
rect 8495 3417 8507 3451
rect 8449 3411 8507 3417
rect 8662 3408 8668 3460
rect 8720 3448 8726 3460
rect 9140 3448 9168 3479
rect 9398 3476 9404 3528
rect 9456 3476 9462 3528
rect 10594 3476 10600 3528
rect 10652 3476 10658 3528
rect 11057 3519 11115 3525
rect 11057 3485 11069 3519
rect 11103 3516 11115 3519
rect 11238 3516 11244 3528
rect 11103 3488 11244 3516
rect 11103 3485 11115 3488
rect 11057 3479 11115 3485
rect 11238 3476 11244 3488
rect 11296 3476 11302 3528
rect 11422 3476 11428 3528
rect 11480 3476 11486 3528
rect 11606 3476 11612 3528
rect 11664 3476 11670 3528
rect 12434 3476 12440 3528
rect 12492 3476 12498 3528
rect 12710 3476 12716 3528
rect 12768 3476 12774 3528
rect 12894 3476 12900 3528
rect 12952 3476 12958 3528
rect 13188 3525 13216 3556
rect 13909 3553 13921 3556
rect 13955 3553 13967 3587
rect 13909 3547 13967 3553
rect 14366 3544 14372 3596
rect 14424 3544 14430 3596
rect 14921 3587 14979 3593
rect 14921 3584 14933 3587
rect 14568 3556 14933 3584
rect 13173 3519 13231 3525
rect 13173 3485 13185 3519
rect 13219 3516 13231 3519
rect 13449 3519 13507 3525
rect 13219 3488 13253 3516
rect 13219 3485 13231 3488
rect 13173 3479 13231 3485
rect 13449 3485 13461 3519
rect 13495 3485 13507 3519
rect 13449 3479 13507 3485
rect 13633 3519 13691 3525
rect 13633 3485 13645 3519
rect 13679 3485 13691 3519
rect 13633 3479 13691 3485
rect 12342 3448 12348 3460
rect 8720 3420 9076 3448
rect 9140 3420 12348 3448
rect 8720 3408 8726 3420
rect 8941 3383 8999 3389
rect 8941 3380 8953 3383
rect 6288 3352 8953 3380
rect 8941 3349 8953 3352
rect 8987 3349 8999 3383
rect 9048 3380 9076 3420
rect 12342 3408 12348 3420
rect 12400 3408 12406 3460
rect 13464 3448 13492 3479
rect 12912 3420 13492 3448
rect 13648 3448 13676 3479
rect 13814 3476 13820 3528
rect 13872 3516 13878 3528
rect 14568 3525 14596 3556
rect 14921 3553 14933 3556
rect 14967 3584 14979 3587
rect 15654 3584 15660 3596
rect 14967 3556 15660 3584
rect 14967 3553 14979 3556
rect 14921 3547 14979 3553
rect 15654 3544 15660 3556
rect 15712 3544 15718 3596
rect 14277 3519 14335 3525
rect 14277 3516 14289 3519
rect 13872 3488 14289 3516
rect 13872 3476 13878 3488
rect 14277 3485 14289 3488
rect 14323 3485 14335 3519
rect 14277 3479 14335 3485
rect 14553 3519 14611 3525
rect 14553 3485 14565 3519
rect 14599 3485 14611 3519
rect 14553 3479 14611 3485
rect 14568 3448 14596 3479
rect 14642 3476 14648 3528
rect 14700 3476 14706 3528
rect 15470 3525 15476 3528
rect 15440 3519 15476 3525
rect 15440 3485 15452 3519
rect 15440 3479 15476 3485
rect 15470 3476 15476 3479
rect 15528 3476 15534 3528
rect 15838 3476 15844 3528
rect 15896 3476 15902 3528
rect 13648 3420 14596 3448
rect 10134 3380 10140 3392
rect 9048 3352 10140 3380
rect 8941 3343 8999 3349
rect 10134 3340 10140 3352
rect 10192 3340 10198 3392
rect 11330 3340 11336 3392
rect 11388 3380 11394 3392
rect 12912 3380 12940 3420
rect 11388 3352 12940 3380
rect 11388 3340 11394 3352
rect 13354 3340 13360 3392
rect 13412 3380 13418 3392
rect 13648 3380 13676 3420
rect 15654 3408 15660 3460
rect 15712 3408 15718 3460
rect 13412 3352 13676 3380
rect 13412 3340 13418 3352
rect 15102 3340 15108 3392
rect 15160 3380 15166 3392
rect 15381 3383 15439 3389
rect 15381 3380 15393 3383
rect 15160 3352 15393 3380
rect 15160 3340 15166 3352
rect 15381 3349 15393 3352
rect 15427 3349 15439 3383
rect 15381 3343 15439 3349
rect 1104 3290 17848 3312
rect 1104 3238 2658 3290
rect 2710 3238 2722 3290
rect 2774 3238 2786 3290
rect 2838 3238 2850 3290
rect 2902 3238 2914 3290
rect 2966 3238 2978 3290
rect 3030 3238 8658 3290
rect 8710 3238 8722 3290
rect 8774 3238 8786 3290
rect 8838 3238 8850 3290
rect 8902 3238 8914 3290
rect 8966 3238 8978 3290
rect 9030 3238 14658 3290
rect 14710 3238 14722 3290
rect 14774 3238 14786 3290
rect 14838 3238 14850 3290
rect 14902 3238 14914 3290
rect 14966 3238 14978 3290
rect 15030 3238 17848 3290
rect 1104 3216 17848 3238
rect 2406 3176 2412 3188
rect 2148 3148 2412 3176
rect 2148 3049 2176 3148
rect 2406 3136 2412 3148
rect 2464 3176 2470 3188
rect 2866 3176 2872 3188
rect 2464 3148 2872 3176
rect 2464 3136 2470 3148
rect 2866 3136 2872 3148
rect 2924 3136 2930 3188
rect 3142 3136 3148 3188
rect 3200 3176 3206 3188
rect 3786 3176 3792 3188
rect 3200 3148 3792 3176
rect 3200 3136 3206 3148
rect 3786 3136 3792 3148
rect 3844 3176 3850 3188
rect 3844 3148 6040 3176
rect 3844 3136 3850 3148
rect 3418 3068 3424 3120
rect 3476 3068 3482 3120
rect 3878 3068 3884 3120
rect 3936 3068 3942 3120
rect 4172 3049 4200 3148
rect 5258 3068 5264 3120
rect 5316 3068 5322 3120
rect 6012 3049 6040 3148
rect 9398 3136 9404 3188
rect 9456 3176 9462 3188
rect 9854 3179 9912 3185
rect 9854 3176 9866 3179
rect 9456 3148 9866 3176
rect 9456 3136 9462 3148
rect 9854 3145 9866 3148
rect 9900 3145 9912 3179
rect 9854 3139 9912 3145
rect 10594 3136 10600 3188
rect 10652 3136 10658 3188
rect 10704 3148 11100 3176
rect 7024 3080 7420 3108
rect 1581 3043 1639 3049
rect 1581 3009 1593 3043
rect 1627 3009 1639 3043
rect 1581 3003 1639 3009
rect 2133 3043 2191 3049
rect 2133 3009 2145 3043
rect 2179 3009 2191 3043
rect 2133 3003 2191 3009
rect 4157 3043 4215 3049
rect 4157 3009 4169 3043
rect 4203 3009 4215 3043
rect 4157 3003 4215 3009
rect 5997 3043 6055 3049
rect 5997 3009 6009 3043
rect 6043 3009 6055 3043
rect 5997 3003 6055 3009
rect 1596 2972 1624 3003
rect 2409 2975 2467 2981
rect 2409 2972 2421 2975
rect 1596 2944 2421 2972
rect 2409 2941 2421 2944
rect 2455 2941 2467 2975
rect 2409 2935 2467 2941
rect 2866 2932 2872 2984
rect 2924 2972 2930 2984
rect 3510 2972 3516 2984
rect 2924 2944 3516 2972
rect 2924 2932 2930 2944
rect 3510 2932 3516 2944
rect 3568 2972 3574 2984
rect 3878 2972 3884 2984
rect 3568 2944 3884 2972
rect 3568 2932 3574 2944
rect 3878 2932 3884 2944
rect 3936 2932 3942 2984
rect 4246 2932 4252 2984
rect 4304 2932 4310 2984
rect 5721 2975 5779 2981
rect 5721 2941 5733 2975
rect 5767 2972 5779 2975
rect 6733 2975 6791 2981
rect 6733 2972 6745 2975
rect 5767 2944 6745 2972
rect 5767 2941 5779 2944
rect 5721 2935 5779 2941
rect 6733 2941 6745 2944
rect 6779 2941 6791 2975
rect 6733 2935 6791 2941
rect 1394 2796 1400 2848
rect 1452 2796 1458 2848
rect 2225 2839 2283 2845
rect 2225 2805 2237 2839
rect 2271 2836 2283 2839
rect 2314 2836 2320 2848
rect 2271 2808 2320 2836
rect 2271 2805 2283 2808
rect 2225 2799 2283 2805
rect 2314 2796 2320 2808
rect 2372 2796 2378 2848
rect 3234 2796 3240 2848
rect 3292 2836 3298 2848
rect 7024 2836 7052 3080
rect 7098 3000 7104 3052
rect 7156 3000 7162 3052
rect 7392 3049 7420 3080
rect 7466 3068 7472 3120
rect 7524 3108 7530 3120
rect 7524 3080 7604 3108
rect 7524 3068 7530 3080
rect 7576 3049 7604 3080
rect 8294 3068 8300 3120
rect 8352 3108 8358 3120
rect 9766 3108 9772 3120
rect 8352 3080 9076 3108
rect 8352 3068 8358 3080
rect 7377 3043 7435 3049
rect 7377 3009 7389 3043
rect 7423 3009 7435 3043
rect 7377 3003 7435 3009
rect 7561 3043 7619 3049
rect 7561 3009 7573 3043
rect 7607 3009 7619 3043
rect 7561 3003 7619 3009
rect 8478 3000 8484 3052
rect 8536 3040 8542 3052
rect 9048 3049 9076 3080
rect 9232 3080 9772 3108
rect 9232 3049 9260 3080
rect 9766 3068 9772 3080
rect 9824 3068 9830 3120
rect 10704 3108 10732 3148
rect 10870 3108 10876 3120
rect 10060 3080 10732 3108
rect 10796 3080 10876 3108
rect 8573 3043 8631 3049
rect 8573 3040 8585 3043
rect 8536 3012 8585 3040
rect 8536 3000 8542 3012
rect 8573 3009 8585 3012
rect 8619 3009 8631 3043
rect 8573 3003 8631 3009
rect 9033 3043 9091 3049
rect 9033 3009 9045 3043
rect 9079 3009 9091 3043
rect 9217 3043 9275 3049
rect 9217 3040 9229 3043
rect 9033 3003 9091 3009
rect 9140 3012 9229 3040
rect 7193 2975 7251 2981
rect 7193 2941 7205 2975
rect 7239 2972 7251 2975
rect 7469 2975 7527 2981
rect 7469 2972 7481 2975
rect 7239 2944 7481 2972
rect 7239 2941 7251 2944
rect 7193 2935 7251 2941
rect 7469 2941 7481 2944
rect 7515 2941 7527 2975
rect 7469 2935 7527 2941
rect 8665 2975 8723 2981
rect 8665 2941 8677 2975
rect 8711 2972 8723 2975
rect 8849 2975 8907 2981
rect 8849 2972 8861 2975
rect 8711 2944 8861 2972
rect 8711 2941 8723 2944
rect 8665 2935 8723 2941
rect 8849 2941 8861 2944
rect 8895 2941 8907 2975
rect 8849 2935 8907 2941
rect 7558 2864 7564 2916
rect 7616 2904 7622 2916
rect 8205 2907 8263 2913
rect 8205 2904 8217 2907
rect 7616 2876 8217 2904
rect 7616 2864 7622 2876
rect 8205 2873 8217 2876
rect 8251 2873 8263 2907
rect 8205 2867 8263 2873
rect 9140 2836 9168 3012
rect 9217 3009 9229 3012
rect 9263 3009 9275 3043
rect 9217 3003 9275 3009
rect 9309 3043 9367 3049
rect 9309 3009 9321 3043
rect 9355 3040 9367 3043
rect 9674 3040 9680 3052
rect 9355 3012 9680 3040
rect 9355 3009 9367 3012
rect 9309 3003 9367 3009
rect 9674 3000 9680 3012
rect 9732 3000 9738 3052
rect 10060 3049 10088 3080
rect 9953 3043 10011 3049
rect 9953 3009 9965 3043
rect 9999 3009 10011 3043
rect 9953 3003 10011 3009
rect 10045 3043 10103 3049
rect 10045 3009 10057 3043
rect 10091 3009 10103 3043
rect 10045 3003 10103 3009
rect 9968 2972 9996 3003
rect 10134 3000 10140 3052
rect 10192 3040 10198 3052
rect 10796 3049 10824 3080
rect 10870 3068 10876 3080
rect 10928 3068 10934 3120
rect 11072 3108 11100 3148
rect 11698 3136 11704 3188
rect 11756 3136 11762 3188
rect 12342 3136 12348 3188
rect 12400 3176 12406 3188
rect 12437 3179 12495 3185
rect 12437 3176 12449 3179
rect 12400 3148 12449 3176
rect 12400 3136 12406 3148
rect 12437 3145 12449 3148
rect 12483 3176 12495 3179
rect 14550 3176 14556 3188
rect 12483 3148 14556 3176
rect 12483 3145 12495 3148
rect 12437 3139 12495 3145
rect 14550 3136 14556 3148
rect 14608 3136 14614 3188
rect 15102 3136 15108 3188
rect 15160 3136 15166 3188
rect 11146 3108 11152 3120
rect 11072 3080 11152 3108
rect 10781 3043 10839 3049
rect 10781 3040 10793 3043
rect 10192 3012 10793 3040
rect 10192 3000 10198 3012
rect 10781 3009 10793 3012
rect 10827 3009 10839 3043
rect 10781 3003 10839 3009
rect 10965 3043 11023 3049
rect 10965 3009 10977 3043
rect 11011 3038 11023 3043
rect 11072 3038 11100 3080
rect 11146 3068 11152 3080
rect 11204 3108 11210 3120
rect 12710 3108 12716 3120
rect 11204 3080 12716 3108
rect 11204 3068 11210 3080
rect 11808 3049 11836 3080
rect 12710 3068 12716 3080
rect 12768 3068 12774 3120
rect 13538 3068 13544 3120
rect 13596 3108 13602 3120
rect 13596 3080 13676 3108
rect 13596 3068 13602 3080
rect 11011 3010 11100 3038
rect 11241 3043 11299 3049
rect 11011 3009 11023 3010
rect 10965 3003 11023 3009
rect 11241 3009 11253 3043
rect 11287 3009 11299 3043
rect 11241 3003 11299 3009
rect 11793 3043 11851 3049
rect 11793 3009 11805 3043
rect 11839 3009 11851 3043
rect 11793 3003 11851 3009
rect 10505 2975 10563 2981
rect 9968 2944 10364 2972
rect 10336 2913 10364 2944
rect 10505 2941 10517 2975
rect 10551 2972 10563 2975
rect 10870 2972 10876 2984
rect 10551 2944 10876 2972
rect 10551 2941 10563 2944
rect 10505 2935 10563 2941
rect 10870 2932 10876 2944
rect 10928 2932 10934 2984
rect 11256 2972 11284 3003
rect 11974 3000 11980 3052
rect 12032 3000 12038 3052
rect 12434 3040 12440 3052
rect 12287 3012 12440 3040
rect 11517 2975 11575 2981
rect 11517 2972 11529 2975
rect 11256 2944 11529 2972
rect 10321 2907 10379 2913
rect 10321 2873 10333 2907
rect 10367 2904 10379 2907
rect 11054 2904 11060 2916
rect 10367 2876 11060 2904
rect 10367 2873 10379 2876
rect 10321 2867 10379 2873
rect 11054 2864 11060 2876
rect 11112 2864 11118 2916
rect 3292 2808 9168 2836
rect 3292 2796 3298 2808
rect 10778 2796 10784 2848
rect 10836 2796 10842 2848
rect 10870 2796 10876 2848
rect 10928 2836 10934 2848
rect 11256 2836 11284 2944
rect 11517 2941 11529 2944
rect 11563 2972 11575 2975
rect 12287 2972 12315 3012
rect 12434 3000 12440 3012
rect 12492 3040 12498 3052
rect 13648 3049 13676 3080
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 12492 3012 13001 3040
rect 12492 3000 12498 3012
rect 12989 3009 13001 3012
rect 13035 3009 13047 3043
rect 12989 3003 13047 3009
rect 13633 3043 13691 3049
rect 13633 3009 13645 3043
rect 13679 3009 13691 3043
rect 13633 3003 13691 3009
rect 13722 3000 13728 3052
rect 13780 3040 13786 3052
rect 14185 3043 14243 3049
rect 14185 3040 14197 3043
rect 13780 3012 14197 3040
rect 13780 3000 13786 3012
rect 14185 3009 14197 3012
rect 14231 3009 14243 3043
rect 14568 3040 14596 3136
rect 15746 3108 15752 3120
rect 15396 3080 15752 3108
rect 15396 3049 15424 3080
rect 15746 3068 15752 3080
rect 15804 3068 15810 3120
rect 15289 3043 15347 3049
rect 15289 3040 15301 3043
rect 14568 3012 15301 3040
rect 14185 3003 14243 3009
rect 15289 3009 15301 3012
rect 15335 3009 15347 3043
rect 15289 3003 15347 3009
rect 15381 3043 15439 3049
rect 15381 3009 15393 3043
rect 15427 3009 15439 3043
rect 15381 3003 15439 3009
rect 15562 3000 15568 3052
rect 15620 3040 15626 3052
rect 15657 3043 15715 3049
rect 15657 3040 15669 3043
rect 15620 3012 15669 3040
rect 15620 3000 15626 3012
rect 15657 3009 15669 3012
rect 15703 3009 15715 3043
rect 15657 3003 15715 3009
rect 12713 2975 12771 2981
rect 12713 2972 12725 2975
rect 11563 2944 12315 2972
rect 12360 2944 12725 2972
rect 11563 2941 11575 2944
rect 11517 2935 11575 2941
rect 11974 2864 11980 2916
rect 12032 2904 12038 2916
rect 12360 2904 12388 2944
rect 12713 2941 12725 2944
rect 12759 2972 12771 2975
rect 12894 2972 12900 2984
rect 12759 2944 12900 2972
rect 12759 2941 12771 2944
rect 12713 2935 12771 2941
rect 12894 2932 12900 2944
rect 12952 2932 12958 2984
rect 14366 2904 14372 2916
rect 12032 2876 12388 2904
rect 12544 2876 14372 2904
rect 12032 2864 12038 2876
rect 10928 2808 11284 2836
rect 10928 2796 10934 2808
rect 12342 2796 12348 2848
rect 12400 2836 12406 2848
rect 12544 2836 12572 2876
rect 14366 2864 14372 2876
rect 14424 2904 14430 2916
rect 15565 2907 15623 2913
rect 15565 2904 15577 2907
rect 14424 2876 15577 2904
rect 14424 2864 14430 2876
rect 15565 2873 15577 2876
rect 15611 2904 15623 2907
rect 15654 2904 15660 2916
rect 15611 2876 15660 2904
rect 15611 2873 15623 2876
rect 15565 2867 15623 2873
rect 15654 2864 15660 2876
rect 15712 2864 15718 2916
rect 12400 2808 12572 2836
rect 12400 2796 12406 2808
rect 12710 2796 12716 2848
rect 12768 2836 12774 2848
rect 12805 2839 12863 2845
rect 12805 2836 12817 2839
rect 12768 2808 12817 2836
rect 12768 2796 12774 2808
rect 12805 2805 12817 2808
rect 12851 2836 12863 2839
rect 13630 2836 13636 2848
rect 12851 2808 13636 2836
rect 12851 2805 12863 2808
rect 12805 2799 12863 2805
rect 13630 2796 13636 2808
rect 13688 2796 13694 2848
rect 1104 2746 17848 2768
rect 1104 2694 1918 2746
rect 1970 2694 1982 2746
rect 2034 2694 2046 2746
rect 2098 2694 2110 2746
rect 2162 2694 2174 2746
rect 2226 2694 2238 2746
rect 2290 2694 7918 2746
rect 7970 2694 7982 2746
rect 8034 2694 8046 2746
rect 8098 2694 8110 2746
rect 8162 2694 8174 2746
rect 8226 2694 8238 2746
rect 8290 2694 13918 2746
rect 13970 2694 13982 2746
rect 14034 2694 14046 2746
rect 14098 2694 14110 2746
rect 14162 2694 14174 2746
rect 14226 2694 14238 2746
rect 14290 2694 17848 2746
rect 1104 2672 17848 2694
rect 1397 2635 1455 2641
rect 1397 2601 1409 2635
rect 1443 2632 1455 2635
rect 1578 2632 1584 2644
rect 1443 2604 1584 2632
rect 1443 2601 1455 2604
rect 1397 2595 1455 2601
rect 1578 2592 1584 2604
rect 1636 2592 1642 2644
rect 3418 2592 3424 2644
rect 3476 2632 3482 2644
rect 3881 2635 3939 2641
rect 3881 2632 3893 2635
rect 3476 2604 3893 2632
rect 3476 2592 3482 2604
rect 3881 2601 3893 2604
rect 3927 2601 3939 2635
rect 3881 2595 3939 2601
rect 5258 2592 5264 2644
rect 5316 2632 5322 2644
rect 5353 2635 5411 2641
rect 5353 2632 5365 2635
rect 5316 2604 5365 2632
rect 5316 2592 5322 2604
rect 5353 2601 5365 2604
rect 5399 2601 5411 2635
rect 5353 2595 5411 2601
rect 9674 2592 9680 2644
rect 9732 2632 9738 2644
rect 11057 2635 11115 2641
rect 11057 2632 11069 2635
rect 9732 2604 11069 2632
rect 9732 2592 9738 2604
rect 11057 2601 11069 2604
rect 11103 2601 11115 2635
rect 11057 2595 11115 2601
rect 13170 2592 13176 2644
rect 13228 2592 13234 2644
rect 12894 2524 12900 2576
rect 12952 2564 12958 2576
rect 12952 2536 13308 2564
rect 12952 2524 12958 2536
rect 3145 2499 3203 2505
rect 3145 2465 3157 2499
rect 3191 2496 3203 2499
rect 3786 2496 3792 2508
rect 3191 2468 3792 2496
rect 3191 2465 3203 2468
rect 3145 2459 3203 2465
rect 3786 2456 3792 2468
rect 3844 2456 3850 2508
rect 9953 2499 10011 2505
rect 9953 2496 9965 2499
rect 6886 2468 9965 2496
rect 3970 2388 3976 2440
rect 4028 2428 4034 2440
rect 5261 2431 5319 2437
rect 5261 2428 5273 2431
rect 4028 2400 5273 2428
rect 4028 2388 4034 2400
rect 5261 2397 5273 2400
rect 5307 2428 5319 2431
rect 6886 2428 6914 2468
rect 9953 2465 9965 2468
rect 9999 2496 10011 2499
rect 12986 2496 12992 2508
rect 9999 2468 12992 2496
rect 9999 2465 10011 2468
rect 9953 2459 10011 2465
rect 12986 2456 12992 2468
rect 13044 2456 13050 2508
rect 5307 2400 6914 2428
rect 5307 2397 5319 2400
rect 5261 2391 5319 2397
rect 9398 2388 9404 2440
rect 9456 2428 9462 2440
rect 9493 2431 9551 2437
rect 9493 2428 9505 2431
rect 9456 2400 9505 2428
rect 9456 2388 9462 2400
rect 9493 2397 9505 2400
rect 9539 2397 9551 2431
rect 9493 2391 9551 2397
rect 11149 2431 11207 2437
rect 11149 2397 11161 2431
rect 11195 2428 11207 2431
rect 11422 2428 11428 2440
rect 11195 2400 11428 2428
rect 11195 2397 11207 2400
rect 11149 2391 11207 2397
rect 11422 2388 11428 2400
rect 11480 2428 11486 2440
rect 12342 2428 12348 2440
rect 11480 2400 12348 2428
rect 11480 2388 11486 2400
rect 12342 2388 12348 2400
rect 12400 2388 12406 2440
rect 12710 2388 12716 2440
rect 12768 2428 12774 2440
rect 13280 2437 13308 2536
rect 13081 2431 13139 2437
rect 13081 2428 13093 2431
rect 12768 2400 13093 2428
rect 12768 2388 12774 2400
rect 13081 2397 13093 2400
rect 13127 2397 13139 2431
rect 13081 2391 13139 2397
rect 13265 2431 13323 2437
rect 13265 2397 13277 2431
rect 13311 2397 13323 2431
rect 13265 2391 13323 2397
rect 2314 2320 2320 2372
rect 2372 2320 2378 2372
rect 2869 2363 2927 2369
rect 2869 2329 2881 2363
rect 2915 2360 2927 2363
rect 7558 2360 7564 2372
rect 2915 2332 7564 2360
rect 2915 2329 2927 2332
rect 2869 2323 2927 2329
rect 7558 2320 7564 2332
rect 7616 2320 7622 2372
rect 1104 2202 17848 2224
rect 1104 2150 2658 2202
rect 2710 2150 2722 2202
rect 2774 2150 2786 2202
rect 2838 2150 2850 2202
rect 2902 2150 2914 2202
rect 2966 2150 2978 2202
rect 3030 2150 8658 2202
rect 8710 2150 8722 2202
rect 8774 2150 8786 2202
rect 8838 2150 8850 2202
rect 8902 2150 8914 2202
rect 8966 2150 8978 2202
rect 9030 2150 14658 2202
rect 14710 2150 14722 2202
rect 14774 2150 14786 2202
rect 14838 2150 14850 2202
rect 14902 2150 14914 2202
rect 14966 2150 14978 2202
rect 15030 2150 17848 2202
rect 1104 2128 17848 2150
<< via1 >>
rect 2658 18470 2710 18522
rect 2722 18470 2774 18522
rect 2786 18470 2838 18522
rect 2850 18470 2902 18522
rect 2914 18470 2966 18522
rect 2978 18470 3030 18522
rect 8658 18470 8710 18522
rect 8722 18470 8774 18522
rect 8786 18470 8838 18522
rect 8850 18470 8902 18522
rect 8914 18470 8966 18522
rect 8978 18470 9030 18522
rect 14658 18470 14710 18522
rect 14722 18470 14774 18522
rect 14786 18470 14838 18522
rect 14850 18470 14902 18522
rect 14914 18470 14966 18522
rect 14978 18470 15030 18522
rect 1216 18368 1268 18420
rect 5724 18368 5776 18420
rect 7012 18368 7064 18420
rect 1124 18232 1176 18284
rect 2228 18232 2280 18284
rect 3332 18232 3384 18284
rect 4436 18232 4488 18284
rect 5540 18232 5592 18284
rect 6644 18300 6696 18352
rect 7104 18300 7156 18352
rect 7932 18232 7984 18284
rect 9128 18232 9180 18284
rect 9956 18232 10008 18284
rect 11060 18275 11112 18284
rect 11060 18241 11069 18275
rect 11069 18241 11103 18275
rect 11103 18241 11112 18275
rect 11060 18232 11112 18241
rect 11152 18275 11204 18284
rect 11152 18241 11161 18275
rect 11161 18241 11195 18275
rect 11195 18241 11204 18275
rect 11152 18232 11204 18241
rect 12164 18232 12216 18284
rect 13268 18232 13320 18284
rect 14372 18232 14424 18284
rect 15476 18232 15528 18284
rect 16580 18232 16632 18284
rect 17684 18232 17736 18284
rect 3516 18164 3568 18216
rect 6368 18207 6420 18216
rect 6368 18173 6377 18207
rect 6377 18173 6411 18207
rect 6411 18173 6420 18207
rect 6368 18164 6420 18173
rect 11980 18164 12032 18216
rect 1584 18071 1636 18080
rect 1584 18037 1593 18071
rect 1593 18037 1627 18071
rect 1627 18037 1636 18071
rect 1584 18028 1636 18037
rect 4896 18028 4948 18080
rect 12164 18096 12216 18148
rect 8484 18071 8536 18080
rect 8484 18037 8493 18071
rect 8493 18037 8527 18071
rect 8527 18037 8536 18071
rect 8484 18028 8536 18037
rect 9956 18028 10008 18080
rect 10048 18071 10100 18080
rect 10048 18037 10057 18071
rect 10057 18037 10091 18071
rect 10091 18037 10100 18071
rect 10048 18028 10100 18037
rect 11060 18028 11112 18080
rect 11796 18028 11848 18080
rect 12440 18071 12492 18080
rect 12440 18037 12449 18071
rect 12449 18037 12483 18071
rect 12483 18037 12492 18071
rect 12440 18028 12492 18037
rect 13268 18028 13320 18080
rect 15476 18028 15528 18080
rect 15568 18071 15620 18080
rect 15568 18037 15577 18071
rect 15577 18037 15611 18071
rect 15611 18037 15620 18071
rect 15568 18028 15620 18037
rect 16028 18028 16080 18080
rect 17224 18028 17276 18080
rect 1918 17926 1970 17978
rect 1982 17926 2034 17978
rect 2046 17926 2098 17978
rect 2110 17926 2162 17978
rect 2174 17926 2226 17978
rect 2238 17926 2290 17978
rect 7918 17926 7970 17978
rect 7982 17926 8034 17978
rect 8046 17926 8098 17978
rect 8110 17926 8162 17978
rect 8174 17926 8226 17978
rect 8238 17926 8290 17978
rect 13918 17926 13970 17978
rect 13982 17926 14034 17978
rect 14046 17926 14098 17978
rect 14110 17926 14162 17978
rect 14174 17926 14226 17978
rect 14238 17926 14290 17978
rect 4068 17688 4120 17740
rect 6368 17688 6420 17740
rect 7012 17731 7064 17740
rect 7012 17697 7021 17731
rect 7021 17697 7055 17731
rect 7055 17697 7064 17731
rect 7012 17688 7064 17697
rect 1584 17552 1636 17604
rect 2228 17552 2280 17604
rect 3240 17552 3292 17604
rect 2504 17484 2556 17536
rect 3884 17527 3936 17536
rect 3884 17493 3893 17527
rect 3893 17493 3927 17527
rect 3927 17493 3936 17527
rect 3884 17484 3936 17493
rect 4436 17527 4488 17536
rect 4436 17493 4445 17527
rect 4445 17493 4479 17527
rect 4479 17493 4488 17527
rect 4436 17484 4488 17493
rect 4896 17595 4948 17604
rect 4896 17561 4905 17595
rect 4905 17561 4939 17595
rect 4939 17561 4948 17595
rect 4896 17552 4948 17561
rect 6460 17552 6512 17604
rect 6644 17595 6696 17604
rect 6644 17561 6653 17595
rect 6653 17561 6687 17595
rect 6687 17561 6696 17595
rect 6644 17552 6696 17561
rect 6552 17484 6604 17536
rect 9772 17731 9824 17740
rect 9772 17697 9781 17731
rect 9781 17697 9815 17731
rect 9815 17697 9824 17731
rect 9772 17688 9824 17697
rect 10048 17731 10100 17740
rect 10048 17697 10057 17731
rect 10057 17697 10091 17731
rect 10091 17697 10100 17731
rect 10048 17688 10100 17697
rect 13544 17688 13596 17740
rect 15568 17688 15620 17740
rect 9128 17663 9180 17672
rect 9128 17629 9137 17663
rect 9137 17629 9171 17663
rect 9171 17629 9180 17663
rect 9128 17620 9180 17629
rect 11060 17552 11112 17604
rect 11428 17552 11480 17604
rect 12164 17595 12216 17604
rect 12164 17561 12173 17595
rect 12173 17561 12207 17595
rect 12207 17561 12216 17595
rect 12164 17552 12216 17561
rect 12624 17552 12676 17604
rect 13452 17552 13504 17604
rect 12256 17484 12308 17536
rect 12348 17484 12400 17536
rect 14556 17620 14608 17672
rect 16764 17620 16816 17672
rect 15660 17552 15712 17604
rect 16488 17552 16540 17604
rect 14280 17484 14332 17536
rect 17040 17484 17092 17536
rect 2658 17382 2710 17434
rect 2722 17382 2774 17434
rect 2786 17382 2838 17434
rect 2850 17382 2902 17434
rect 2914 17382 2966 17434
rect 2978 17382 3030 17434
rect 8658 17382 8710 17434
rect 8722 17382 8774 17434
rect 8786 17382 8838 17434
rect 8850 17382 8902 17434
rect 8914 17382 8966 17434
rect 8978 17382 9030 17434
rect 14658 17382 14710 17434
rect 14722 17382 14774 17434
rect 14786 17382 14838 17434
rect 14850 17382 14902 17434
rect 14914 17382 14966 17434
rect 14978 17382 15030 17434
rect 1308 17280 1360 17332
rect 2228 17323 2280 17332
rect 2228 17289 2237 17323
rect 2237 17289 2271 17323
rect 2271 17289 2280 17323
rect 2228 17280 2280 17289
rect 3516 17323 3568 17332
rect 3516 17289 3525 17323
rect 3525 17289 3559 17323
rect 3559 17289 3568 17323
rect 3516 17280 3568 17289
rect 6460 17323 6512 17332
rect 6460 17289 6469 17323
rect 6469 17289 6503 17323
rect 6503 17289 6512 17323
rect 6460 17280 6512 17289
rect 7104 17323 7156 17332
rect 7104 17289 7113 17323
rect 7113 17289 7147 17323
rect 7147 17289 7156 17323
rect 7104 17280 7156 17289
rect 9128 17280 9180 17332
rect 4436 17212 4488 17264
rect 8484 17212 8536 17264
rect 9220 17212 9272 17264
rect 2504 17144 2556 17196
rect 6552 17187 6604 17196
rect 6552 17153 6561 17187
rect 6561 17153 6595 17187
rect 6595 17153 6604 17187
rect 11152 17280 11204 17332
rect 12624 17280 12676 17332
rect 15660 17323 15712 17332
rect 15660 17289 15669 17323
rect 15669 17289 15703 17323
rect 15703 17289 15712 17323
rect 15660 17280 15712 17289
rect 6552 17144 6604 17153
rect 12348 17144 12400 17196
rect 13544 17212 13596 17264
rect 14280 17212 14332 17264
rect 14556 17144 14608 17196
rect 16764 17144 16816 17196
rect 3056 17076 3108 17128
rect 4252 17076 4304 17128
rect 3976 16940 4028 16992
rect 9864 17076 9916 17128
rect 12072 17076 12124 17128
rect 13268 17119 13320 17128
rect 13268 17085 13277 17119
rect 13277 17085 13311 17119
rect 13311 17085 13320 17119
rect 13268 17076 13320 17085
rect 16856 17076 16908 17128
rect 11152 16940 11204 16992
rect 1918 16838 1970 16890
rect 1982 16838 2034 16890
rect 2046 16838 2098 16890
rect 2110 16838 2162 16890
rect 2174 16838 2226 16890
rect 2238 16838 2290 16890
rect 7918 16838 7970 16890
rect 7982 16838 8034 16890
rect 8046 16838 8098 16890
rect 8110 16838 8162 16890
rect 8174 16838 8226 16890
rect 8238 16838 8290 16890
rect 13918 16838 13970 16890
rect 13982 16838 14034 16890
rect 14046 16838 14098 16890
rect 14110 16838 14162 16890
rect 14174 16838 14226 16890
rect 14238 16838 14290 16890
rect 4344 16736 4396 16788
rect 9220 16736 9272 16788
rect 9956 16736 10008 16788
rect 3332 16600 3384 16652
rect 1400 16532 1452 16584
rect 4068 16575 4120 16584
rect 4068 16541 4077 16575
rect 4077 16541 4111 16575
rect 4111 16541 4120 16575
rect 4068 16532 4120 16541
rect 13912 16668 13964 16720
rect 5816 16600 5868 16652
rect 9128 16600 9180 16652
rect 9864 16643 9916 16652
rect 9864 16609 9873 16643
rect 9873 16609 9907 16643
rect 9907 16609 9916 16643
rect 9864 16600 9916 16609
rect 10140 16600 10192 16652
rect 13544 16600 13596 16652
rect 16028 16643 16080 16652
rect 16028 16609 16037 16643
rect 16037 16609 16071 16643
rect 16071 16609 16080 16643
rect 16028 16600 16080 16609
rect 848 16396 900 16448
rect 4160 16396 4212 16448
rect 12992 16575 13044 16584
rect 12992 16541 13001 16575
rect 13001 16541 13035 16575
rect 13035 16541 13044 16575
rect 12992 16532 13044 16541
rect 13912 16532 13964 16584
rect 11152 16464 11204 16516
rect 12440 16464 12492 16516
rect 15568 16575 15620 16584
rect 15568 16541 15577 16575
rect 15577 16541 15611 16575
rect 15611 16541 15620 16575
rect 15568 16532 15620 16541
rect 6552 16396 6604 16448
rect 12808 16439 12860 16448
rect 12808 16405 12817 16439
rect 12817 16405 12851 16439
rect 12851 16405 12860 16439
rect 12808 16396 12860 16405
rect 13452 16396 13504 16448
rect 15108 16396 15160 16448
rect 17040 16464 17092 16516
rect 15568 16396 15620 16448
rect 15844 16396 15896 16448
rect 2658 16294 2710 16346
rect 2722 16294 2774 16346
rect 2786 16294 2838 16346
rect 2850 16294 2902 16346
rect 2914 16294 2966 16346
rect 2978 16294 3030 16346
rect 8658 16294 8710 16346
rect 8722 16294 8774 16346
rect 8786 16294 8838 16346
rect 8850 16294 8902 16346
rect 8914 16294 8966 16346
rect 8978 16294 9030 16346
rect 14658 16294 14710 16346
rect 14722 16294 14774 16346
rect 14786 16294 14838 16346
rect 14850 16294 14902 16346
rect 14914 16294 14966 16346
rect 14978 16294 15030 16346
rect 3056 16192 3108 16244
rect 4068 16192 4120 16244
rect 5816 16235 5868 16244
rect 5816 16201 5825 16235
rect 5825 16201 5859 16235
rect 5859 16201 5868 16235
rect 5816 16192 5868 16201
rect 7288 16192 7340 16244
rect 7840 16192 7892 16244
rect 12348 16192 12400 16244
rect 3884 16124 3936 16176
rect 4344 16167 4396 16176
rect 4344 16133 4353 16167
rect 4353 16133 4387 16167
rect 4387 16133 4396 16167
rect 4344 16124 4396 16133
rect 1584 16099 1636 16108
rect 1584 16065 1593 16099
rect 1593 16065 1627 16099
rect 1627 16065 1636 16099
rect 1584 16056 1636 16065
rect 2504 16056 2556 16108
rect 3148 15988 3200 16040
rect 3976 15988 4028 16040
rect 6552 16099 6604 16108
rect 6552 16065 6561 16099
rect 6561 16065 6595 16099
rect 6595 16065 6604 16099
rect 6552 16056 6604 16065
rect 7104 16056 7156 16108
rect 7288 16099 7340 16108
rect 7288 16065 7297 16099
rect 7297 16065 7331 16099
rect 7331 16065 7340 16099
rect 7288 16056 7340 16065
rect 9588 16124 9640 16176
rect 8852 16099 8904 16108
rect 8852 16065 8861 16099
rect 8861 16065 8895 16099
rect 8895 16065 8904 16099
rect 8852 16056 8904 16065
rect 12256 16099 12308 16108
rect 12256 16065 12265 16099
rect 12265 16065 12299 16099
rect 12299 16065 12308 16099
rect 12256 16056 12308 16065
rect 12532 16124 12584 16176
rect 14004 16192 14056 16244
rect 14464 16192 14516 16244
rect 14832 16192 14884 16244
rect 15108 16192 15160 16244
rect 15568 16124 15620 16176
rect 12808 16099 12860 16108
rect 12808 16065 12817 16099
rect 12817 16065 12851 16099
rect 12851 16065 12860 16099
rect 12808 16056 12860 16065
rect 12992 16056 13044 16108
rect 7748 15920 7800 15972
rect 13084 15988 13136 16040
rect 13360 15988 13412 16040
rect 13912 16099 13964 16108
rect 13912 16065 13921 16099
rect 13921 16065 13955 16099
rect 13955 16065 13964 16099
rect 13912 16056 13964 16065
rect 14004 16099 14056 16108
rect 14004 16065 14013 16099
rect 14013 16065 14047 16099
rect 14047 16065 14056 16099
rect 14004 16056 14056 16065
rect 13820 15920 13872 15972
rect 14832 16099 14884 16108
rect 14832 16065 14841 16099
rect 14841 16065 14875 16099
rect 14875 16065 14884 16099
rect 14832 16056 14884 16065
rect 14924 16099 14976 16108
rect 14924 16065 14933 16099
rect 14933 16065 14967 16099
rect 14967 16065 14976 16099
rect 14924 16056 14976 16065
rect 16488 16124 16540 16176
rect 15016 15988 15068 16040
rect 15844 16099 15896 16108
rect 15844 16065 15853 16099
rect 15853 16065 15887 16099
rect 15887 16065 15896 16099
rect 15844 16056 15896 16065
rect 16764 16056 16816 16108
rect 15292 15988 15344 16040
rect 14832 15920 14884 15972
rect 848 15852 900 15904
rect 2320 15852 2372 15904
rect 9588 15852 9640 15904
rect 11704 15852 11756 15904
rect 12164 15852 12216 15904
rect 13360 15852 13412 15904
rect 16948 15895 17000 15904
rect 16948 15861 16957 15895
rect 16957 15861 16991 15895
rect 16991 15861 17000 15895
rect 16948 15852 17000 15861
rect 1918 15750 1970 15802
rect 1982 15750 2034 15802
rect 2046 15750 2098 15802
rect 2110 15750 2162 15802
rect 2174 15750 2226 15802
rect 2238 15750 2290 15802
rect 7918 15750 7970 15802
rect 7982 15750 8034 15802
rect 8046 15750 8098 15802
rect 8110 15750 8162 15802
rect 8174 15750 8226 15802
rect 8238 15750 8290 15802
rect 13918 15750 13970 15802
rect 13982 15750 14034 15802
rect 14046 15750 14098 15802
rect 14110 15750 14162 15802
rect 14174 15750 14226 15802
rect 14238 15750 14290 15802
rect 1400 15691 1452 15700
rect 1400 15657 1409 15691
rect 1409 15657 1443 15691
rect 1443 15657 1452 15691
rect 1400 15648 1452 15657
rect 3332 15691 3384 15700
rect 3332 15657 3341 15691
rect 3341 15657 3375 15691
rect 3375 15657 3384 15691
rect 3332 15648 3384 15657
rect 3148 15487 3200 15496
rect 3148 15453 3157 15487
rect 3157 15453 3191 15487
rect 3191 15453 3200 15487
rect 3148 15444 3200 15453
rect 4252 15555 4304 15564
rect 4252 15521 4261 15555
rect 4261 15521 4295 15555
rect 4295 15521 4304 15555
rect 4252 15512 4304 15521
rect 8852 15648 8904 15700
rect 11704 15648 11756 15700
rect 13636 15648 13688 15700
rect 7012 15580 7064 15632
rect 7472 15512 7524 15564
rect 9220 15512 9272 15564
rect 11612 15580 11664 15632
rect 2320 15376 2372 15428
rect 7656 15487 7708 15496
rect 7656 15453 7679 15487
rect 7679 15453 7708 15487
rect 7656 15444 7708 15453
rect 7012 15419 7064 15428
rect 7012 15385 7021 15419
rect 7021 15385 7055 15419
rect 7055 15385 7064 15419
rect 7012 15376 7064 15385
rect 9128 15487 9180 15496
rect 9128 15453 9134 15487
rect 9134 15453 9168 15487
rect 9168 15453 9180 15487
rect 12624 15580 12676 15632
rect 9128 15444 9180 15453
rect 9588 15487 9640 15496
rect 9588 15453 9597 15487
rect 9597 15453 9631 15487
rect 9631 15453 9640 15487
rect 9588 15444 9640 15453
rect 9956 15487 10008 15496
rect 9956 15453 9965 15487
rect 9965 15453 9999 15487
rect 9999 15453 10008 15487
rect 9956 15444 10008 15453
rect 10416 15444 10468 15496
rect 14096 15512 14148 15564
rect 14924 15580 14976 15632
rect 15108 15580 15160 15632
rect 14556 15512 14608 15564
rect 11612 15487 11664 15496
rect 11612 15453 11621 15487
rect 11621 15453 11655 15487
rect 11655 15453 11664 15487
rect 11612 15444 11664 15453
rect 11244 15376 11296 15428
rect 6920 15308 6972 15360
rect 8300 15308 8352 15360
rect 9220 15308 9272 15360
rect 10416 15351 10468 15360
rect 10416 15317 10425 15351
rect 10425 15317 10459 15351
rect 10459 15317 10468 15351
rect 10416 15308 10468 15317
rect 10508 15351 10560 15360
rect 10508 15317 10517 15351
rect 10517 15317 10551 15351
rect 10551 15317 10560 15351
rect 10508 15308 10560 15317
rect 12348 15487 12400 15496
rect 12348 15453 12357 15487
rect 12357 15453 12391 15487
rect 12391 15453 12400 15487
rect 12348 15444 12400 15453
rect 12440 15487 12492 15496
rect 12440 15453 12449 15487
rect 12449 15453 12483 15487
rect 12483 15453 12492 15487
rect 12440 15444 12492 15453
rect 12624 15444 12676 15496
rect 12716 15487 12768 15496
rect 12716 15453 12725 15487
rect 12725 15453 12759 15487
rect 12759 15453 12768 15487
rect 12716 15444 12768 15453
rect 13360 15487 13412 15496
rect 13360 15453 13369 15487
rect 13369 15453 13403 15487
rect 13403 15453 13412 15487
rect 13360 15444 13412 15453
rect 13176 15419 13228 15428
rect 13176 15385 13185 15419
rect 13185 15385 13219 15419
rect 13219 15385 13228 15419
rect 13176 15376 13228 15385
rect 13820 15376 13872 15428
rect 14832 15487 14884 15496
rect 14832 15453 14841 15487
rect 14841 15453 14875 15487
rect 14875 15453 14884 15487
rect 14832 15444 14884 15453
rect 14924 15487 14976 15496
rect 14924 15453 14933 15487
rect 14933 15453 14967 15487
rect 14967 15453 14976 15487
rect 14924 15444 14976 15453
rect 15108 15487 15160 15496
rect 15108 15453 15117 15487
rect 15117 15453 15151 15487
rect 15151 15453 15160 15487
rect 15108 15444 15160 15453
rect 17224 15555 17276 15564
rect 17224 15521 17233 15555
rect 17233 15521 17267 15555
rect 17267 15521 17276 15555
rect 17224 15512 17276 15521
rect 17500 15487 17552 15496
rect 17500 15453 17509 15487
rect 17509 15453 17543 15487
rect 17543 15453 17552 15487
rect 17500 15444 17552 15453
rect 12532 15308 12584 15360
rect 12716 15308 12768 15360
rect 14924 15308 14976 15360
rect 15660 15376 15712 15428
rect 16948 15376 17000 15428
rect 2658 15206 2710 15258
rect 2722 15206 2774 15258
rect 2786 15206 2838 15258
rect 2850 15206 2902 15258
rect 2914 15206 2966 15258
rect 2978 15206 3030 15258
rect 8658 15206 8710 15258
rect 8722 15206 8774 15258
rect 8786 15206 8838 15258
rect 8850 15206 8902 15258
rect 8914 15206 8966 15258
rect 8978 15206 9030 15258
rect 14658 15206 14710 15258
rect 14722 15206 14774 15258
rect 14786 15206 14838 15258
rect 14850 15206 14902 15258
rect 14914 15206 14966 15258
rect 14978 15206 15030 15258
rect 1584 15104 1636 15156
rect 4252 15147 4304 15156
rect 4252 15113 4261 15147
rect 4261 15113 4295 15147
rect 4295 15113 4304 15147
rect 4252 15104 4304 15113
rect 7840 15104 7892 15156
rect 2412 15036 2464 15088
rect 6920 15079 6972 15088
rect 6920 15045 6929 15079
rect 6929 15045 6963 15079
rect 6963 15045 6972 15079
rect 6920 15036 6972 15045
rect 7748 15036 7800 15088
rect 9588 15104 9640 15156
rect 10416 15104 10468 15156
rect 12532 15104 12584 15156
rect 13176 15104 13228 15156
rect 14372 15104 14424 15156
rect 15292 15104 15344 15156
rect 4068 14968 4120 15020
rect 7472 15011 7524 15020
rect 7472 14977 7481 15011
rect 7481 14977 7515 15011
rect 7515 14977 7524 15011
rect 7472 14968 7524 14977
rect 7656 15011 7708 15020
rect 7656 14977 7665 15011
rect 7665 14977 7699 15011
rect 7699 14977 7708 15011
rect 7656 14968 7708 14977
rect 9128 15036 9180 15088
rect 8300 14968 8352 15020
rect 10508 15036 10560 15088
rect 11152 14968 11204 15020
rect 12164 15011 12216 15020
rect 12164 14977 12173 15011
rect 12173 14977 12207 15011
rect 12207 14977 12216 15011
rect 12164 14968 12216 14977
rect 13636 15036 13688 15088
rect 14464 15036 14516 15088
rect 2872 14943 2924 14952
rect 2872 14909 2881 14943
rect 2881 14909 2915 14943
rect 2915 14909 2924 14943
rect 2872 14900 2924 14909
rect 3148 14943 3200 14952
rect 3148 14909 3157 14943
rect 3157 14909 3191 14943
rect 3191 14909 3200 14943
rect 3148 14900 3200 14909
rect 4436 14943 4488 14952
rect 4436 14909 4445 14943
rect 4445 14909 4479 14943
rect 4479 14909 4488 14943
rect 4436 14900 4488 14909
rect 4620 14943 4672 14952
rect 4620 14909 4629 14943
rect 4629 14909 4663 14943
rect 4663 14909 4672 14943
rect 4620 14900 4672 14909
rect 5356 14900 5408 14952
rect 9956 14900 10008 14952
rect 7012 14832 7064 14884
rect 10876 14900 10928 14952
rect 12716 15011 12768 15020
rect 12716 14977 12725 15011
rect 12725 14977 12759 15011
rect 12759 14977 12768 15011
rect 12716 14968 12768 14977
rect 12808 14968 12860 15020
rect 13176 14900 13228 14952
rect 13360 14900 13412 14952
rect 14556 15011 14608 15020
rect 14556 14977 14565 15011
rect 14565 14977 14599 15011
rect 14599 14977 14608 15011
rect 14556 14968 14608 14977
rect 13084 14832 13136 14884
rect 14096 14875 14148 14884
rect 14096 14841 14105 14875
rect 14105 14841 14139 14875
rect 14139 14841 14148 14875
rect 14096 14832 14148 14841
rect 14648 14943 14700 14952
rect 14648 14909 14657 14943
rect 14657 14909 14691 14943
rect 14691 14909 14700 14943
rect 14648 14900 14700 14909
rect 15108 14900 15160 14952
rect 15384 14968 15436 15020
rect 15660 15011 15712 15020
rect 15660 14977 15669 15011
rect 15669 14977 15703 15011
rect 15703 14977 15712 15011
rect 15660 14968 15712 14977
rect 16764 14968 16816 15020
rect 15936 14832 15988 14884
rect 6092 14764 6144 14816
rect 8668 14807 8720 14816
rect 8668 14773 8677 14807
rect 8677 14773 8711 14807
rect 8711 14773 8720 14807
rect 8668 14764 8720 14773
rect 8760 14764 8812 14816
rect 11060 14764 11112 14816
rect 12808 14764 12860 14816
rect 13728 14764 13780 14816
rect 14648 14764 14700 14816
rect 15108 14764 15160 14816
rect 15292 14764 15344 14816
rect 16028 14807 16080 14816
rect 16028 14773 16037 14807
rect 16037 14773 16071 14807
rect 16071 14773 16080 14807
rect 16028 14764 16080 14773
rect 16672 14764 16724 14816
rect 1918 14662 1970 14714
rect 1982 14662 2034 14714
rect 2046 14662 2098 14714
rect 2110 14662 2162 14714
rect 2174 14662 2226 14714
rect 2238 14662 2290 14714
rect 7918 14662 7970 14714
rect 7982 14662 8034 14714
rect 8046 14662 8098 14714
rect 8110 14662 8162 14714
rect 8174 14662 8226 14714
rect 8238 14662 8290 14714
rect 13918 14662 13970 14714
rect 13982 14662 14034 14714
rect 14046 14662 14098 14714
rect 14110 14662 14162 14714
rect 14174 14662 14226 14714
rect 14238 14662 14290 14714
rect 2412 14603 2464 14612
rect 2412 14569 2421 14603
rect 2421 14569 2455 14603
rect 2455 14569 2464 14603
rect 2412 14560 2464 14569
rect 2872 14560 2924 14612
rect 4344 14560 4396 14612
rect 5356 14560 5408 14612
rect 8668 14560 8720 14612
rect 9220 14560 9272 14612
rect 10876 14603 10928 14612
rect 10876 14569 10885 14603
rect 10885 14569 10919 14603
rect 10919 14569 10928 14603
rect 10876 14560 10928 14569
rect 11060 14603 11112 14612
rect 11060 14569 11069 14603
rect 11069 14569 11103 14603
rect 11103 14569 11112 14603
rect 11060 14560 11112 14569
rect 11244 14560 11296 14612
rect 12256 14560 12308 14612
rect 13360 14560 13412 14612
rect 1400 14356 1452 14408
rect 2504 14399 2556 14408
rect 2504 14365 2513 14399
rect 2513 14365 2547 14399
rect 2547 14365 2556 14399
rect 2504 14356 2556 14365
rect 4160 14399 4212 14408
rect 4160 14365 4169 14399
rect 4169 14365 4203 14399
rect 4203 14365 4212 14399
rect 4160 14356 4212 14365
rect 4988 14399 5040 14408
rect 4068 14288 4120 14340
rect 4436 14331 4488 14340
rect 848 14220 900 14272
rect 4160 14220 4212 14272
rect 4436 14297 4463 14331
rect 4463 14297 4488 14331
rect 4988 14365 4997 14399
rect 4997 14365 5031 14399
rect 5031 14365 5040 14399
rect 4988 14356 5040 14365
rect 5356 14399 5408 14408
rect 5356 14365 5365 14399
rect 5365 14365 5399 14399
rect 5399 14365 5408 14399
rect 5356 14356 5408 14365
rect 6092 14492 6144 14544
rect 4436 14288 4488 14297
rect 4620 14331 4672 14340
rect 4620 14297 4629 14331
rect 4629 14297 4663 14331
rect 4663 14297 4672 14331
rect 4620 14288 4672 14297
rect 6092 14399 6144 14408
rect 6092 14365 6101 14399
rect 6101 14365 6135 14399
rect 6135 14365 6144 14399
rect 6092 14356 6144 14365
rect 9864 14424 9916 14476
rect 13820 14424 13872 14476
rect 6828 14356 6880 14408
rect 8760 14356 8812 14408
rect 9772 14356 9824 14408
rect 6920 14288 6972 14340
rect 10692 14356 10744 14408
rect 10876 14356 10928 14408
rect 11152 14399 11204 14408
rect 11152 14365 11161 14399
rect 11161 14365 11195 14399
rect 11195 14365 11204 14399
rect 11152 14356 11204 14365
rect 13544 14356 13596 14408
rect 17500 14424 17552 14476
rect 15476 14288 15528 14340
rect 16672 14288 16724 14340
rect 17408 14263 17460 14272
rect 17408 14229 17417 14263
rect 17417 14229 17451 14263
rect 17451 14229 17460 14263
rect 17408 14220 17460 14229
rect 2658 14118 2710 14170
rect 2722 14118 2774 14170
rect 2786 14118 2838 14170
rect 2850 14118 2902 14170
rect 2914 14118 2966 14170
rect 2978 14118 3030 14170
rect 8658 14118 8710 14170
rect 8722 14118 8774 14170
rect 8786 14118 8838 14170
rect 8850 14118 8902 14170
rect 8914 14118 8966 14170
rect 8978 14118 9030 14170
rect 14658 14118 14710 14170
rect 14722 14118 14774 14170
rect 14786 14118 14838 14170
rect 14850 14118 14902 14170
rect 14914 14118 14966 14170
rect 14978 14118 15030 14170
rect 1400 14059 1452 14068
rect 1400 14025 1409 14059
rect 1409 14025 1443 14059
rect 1443 14025 1452 14059
rect 1400 14016 1452 14025
rect 9772 14059 9824 14068
rect 9772 14025 9781 14059
rect 9781 14025 9815 14059
rect 9815 14025 9824 14059
rect 9772 14016 9824 14025
rect 2320 13948 2372 14000
rect 6920 13880 6972 13932
rect 9496 13880 9548 13932
rect 2872 13855 2924 13864
rect 2872 13821 2881 13855
rect 2881 13821 2915 13855
rect 2915 13821 2924 13855
rect 2872 13812 2924 13821
rect 3148 13855 3200 13864
rect 3148 13821 3157 13855
rect 3157 13821 3191 13855
rect 3191 13821 3200 13855
rect 3148 13812 3200 13821
rect 6828 13855 6880 13864
rect 6828 13821 6837 13855
rect 6837 13821 6871 13855
rect 6871 13821 6880 13855
rect 6828 13812 6880 13821
rect 9312 13855 9364 13864
rect 9312 13821 9321 13855
rect 9321 13821 9355 13855
rect 9355 13821 9364 13855
rect 9312 13812 9364 13821
rect 9864 13923 9916 13932
rect 9864 13889 9873 13923
rect 9873 13889 9907 13923
rect 9907 13889 9916 13923
rect 9864 13880 9916 13889
rect 10968 14016 11020 14068
rect 11060 14016 11112 14068
rect 11612 14016 11664 14068
rect 13268 14016 13320 14068
rect 13452 14059 13504 14068
rect 13452 14025 13461 14059
rect 13461 14025 13495 14059
rect 13495 14025 13504 14059
rect 13452 14016 13504 14025
rect 14372 14016 14424 14068
rect 14648 13948 14700 14000
rect 9588 13744 9640 13796
rect 10692 13855 10744 13864
rect 10692 13821 10701 13855
rect 10701 13821 10735 13855
rect 10735 13821 10744 13855
rect 10692 13812 10744 13821
rect 11244 13923 11296 13932
rect 11244 13889 11253 13923
rect 11253 13889 11287 13923
rect 11287 13889 11296 13923
rect 11244 13880 11296 13889
rect 13084 13923 13136 13932
rect 13084 13889 13093 13923
rect 13093 13889 13127 13923
rect 13127 13889 13136 13923
rect 13084 13880 13136 13889
rect 13360 13923 13412 13932
rect 13360 13889 13369 13923
rect 13369 13889 13403 13923
rect 13403 13889 13412 13923
rect 13360 13880 13412 13889
rect 13728 13880 13780 13932
rect 11336 13744 11388 13796
rect 12348 13744 12400 13796
rect 12532 13744 12584 13796
rect 13912 13812 13964 13864
rect 15752 14016 15804 14068
rect 15292 13948 15344 14000
rect 15108 13880 15160 13932
rect 14464 13744 14516 13796
rect 15384 13880 15436 13932
rect 16028 13880 16080 13932
rect 16856 13880 16908 13932
rect 16580 13812 16632 13864
rect 15660 13744 15712 13796
rect 6368 13676 6420 13728
rect 8484 13676 8536 13728
rect 14924 13719 14976 13728
rect 14924 13685 14933 13719
rect 14933 13685 14967 13719
rect 14967 13685 14976 13719
rect 14924 13676 14976 13685
rect 15384 13719 15436 13728
rect 15384 13685 15393 13719
rect 15393 13685 15427 13719
rect 15427 13685 15436 13719
rect 15384 13676 15436 13685
rect 15476 13719 15528 13728
rect 15476 13685 15485 13719
rect 15485 13685 15519 13719
rect 15519 13685 15528 13719
rect 15476 13676 15528 13685
rect 17408 13676 17460 13728
rect 1918 13574 1970 13626
rect 1982 13574 2034 13626
rect 2046 13574 2098 13626
rect 2110 13574 2162 13626
rect 2174 13574 2226 13626
rect 2238 13574 2290 13626
rect 7918 13574 7970 13626
rect 7982 13574 8034 13626
rect 8046 13574 8098 13626
rect 8110 13574 8162 13626
rect 8174 13574 8226 13626
rect 8238 13574 8290 13626
rect 13918 13574 13970 13626
rect 13982 13574 14034 13626
rect 14046 13574 14098 13626
rect 14110 13574 14162 13626
rect 14174 13574 14226 13626
rect 14238 13574 14290 13626
rect 2320 13515 2372 13524
rect 2320 13481 2329 13515
rect 2329 13481 2363 13515
rect 2363 13481 2372 13515
rect 2320 13472 2372 13481
rect 2872 13472 2924 13524
rect 5264 13472 5316 13524
rect 7656 13472 7708 13524
rect 11152 13515 11204 13524
rect 11152 13481 11161 13515
rect 11161 13481 11195 13515
rect 11195 13481 11204 13515
rect 11152 13472 11204 13481
rect 13268 13472 13320 13524
rect 13912 13472 13964 13524
rect 5356 13379 5408 13388
rect 1400 13268 1452 13320
rect 2504 13268 2556 13320
rect 3516 13268 3568 13320
rect 5356 13345 5365 13379
rect 5365 13345 5399 13379
rect 5399 13345 5408 13379
rect 5356 13336 5408 13345
rect 5264 13311 5316 13320
rect 5264 13277 5266 13311
rect 5266 13277 5300 13311
rect 5300 13277 5316 13311
rect 5264 13268 5316 13277
rect 5632 13311 5684 13320
rect 5632 13277 5641 13311
rect 5641 13277 5675 13311
rect 5675 13277 5684 13311
rect 5632 13268 5684 13277
rect 6368 13311 6420 13320
rect 6368 13277 6377 13311
rect 6377 13277 6411 13311
rect 6411 13277 6420 13311
rect 6368 13268 6420 13277
rect 7748 13336 7800 13388
rect 7104 13268 7156 13320
rect 7564 13311 7616 13320
rect 7564 13277 7573 13311
rect 7573 13277 7607 13311
rect 7607 13277 7616 13311
rect 7564 13268 7616 13277
rect 13820 13404 13872 13456
rect 14648 13404 14700 13456
rect 9496 13336 9548 13388
rect 11060 13336 11112 13388
rect 11980 13336 12032 13388
rect 12808 13336 12860 13388
rect 14924 13336 14976 13388
rect 10140 13268 10192 13320
rect 11336 13311 11388 13320
rect 11336 13277 11345 13311
rect 11345 13277 11379 13311
rect 11379 13277 11388 13311
rect 11336 13268 11388 13277
rect 12164 13268 12216 13320
rect 13544 13311 13596 13320
rect 13544 13277 13553 13311
rect 13553 13277 13587 13311
rect 13587 13277 13596 13311
rect 13544 13268 13596 13277
rect 14464 13268 14516 13320
rect 14740 13311 14792 13320
rect 14740 13277 14749 13311
rect 14749 13277 14783 13311
rect 14783 13277 14792 13311
rect 14740 13268 14792 13277
rect 9680 13200 9732 13252
rect 14280 13200 14332 13252
rect 15384 13311 15436 13320
rect 15384 13277 15393 13311
rect 15393 13277 15427 13311
rect 15427 13277 15436 13311
rect 15384 13268 15436 13277
rect 16396 13379 16448 13388
rect 16396 13345 16405 13379
rect 16405 13345 16439 13379
rect 16439 13345 16448 13379
rect 16396 13336 16448 13345
rect 17408 13336 17460 13388
rect 16580 13268 16632 13320
rect 16764 13311 16816 13320
rect 16764 13277 16773 13311
rect 16773 13277 16807 13311
rect 16807 13277 16816 13311
rect 16764 13268 16816 13277
rect 16856 13311 16908 13320
rect 16856 13277 16865 13311
rect 16865 13277 16899 13311
rect 16899 13277 16908 13311
rect 16856 13268 16908 13277
rect 848 13132 900 13184
rect 4988 13132 5040 13184
rect 6368 13132 6420 13184
rect 12072 13132 12124 13184
rect 12716 13132 12768 13184
rect 13544 13132 13596 13184
rect 13728 13132 13780 13184
rect 14464 13132 14516 13184
rect 14740 13132 14792 13184
rect 16212 13132 16264 13184
rect 2658 13030 2710 13082
rect 2722 13030 2774 13082
rect 2786 13030 2838 13082
rect 2850 13030 2902 13082
rect 2914 13030 2966 13082
rect 2978 13030 3030 13082
rect 8658 13030 8710 13082
rect 8722 13030 8774 13082
rect 8786 13030 8838 13082
rect 8850 13030 8902 13082
rect 8914 13030 8966 13082
rect 8978 13030 9030 13082
rect 14658 13030 14710 13082
rect 14722 13030 14774 13082
rect 14786 13030 14838 13082
rect 14850 13030 14902 13082
rect 14914 13030 14966 13082
rect 14978 13030 15030 13082
rect 1400 12971 1452 12980
rect 1400 12937 1409 12971
rect 1409 12937 1443 12971
rect 1443 12937 1452 12971
rect 1400 12928 1452 12937
rect 3516 12971 3568 12980
rect 3516 12937 3525 12971
rect 3525 12937 3559 12971
rect 3559 12937 3568 12971
rect 3516 12928 3568 12937
rect 5356 12928 5408 12980
rect 2320 12860 2372 12912
rect 3424 12835 3476 12844
rect 3424 12801 3433 12835
rect 3433 12801 3467 12835
rect 3467 12801 3476 12835
rect 3424 12792 3476 12801
rect 4712 12835 4764 12844
rect 4712 12801 4751 12835
rect 4751 12801 4764 12835
rect 4712 12792 4764 12801
rect 3608 12656 3660 12708
rect 4252 12656 4304 12708
rect 4988 12767 5040 12776
rect 4988 12733 4997 12767
rect 4997 12733 5031 12767
rect 5031 12733 5040 12767
rect 4988 12724 5040 12733
rect 5172 12792 5224 12844
rect 5356 12835 5408 12844
rect 5356 12801 5365 12835
rect 5365 12801 5399 12835
rect 5399 12801 5408 12835
rect 5356 12792 5408 12801
rect 7564 12928 7616 12980
rect 9588 12928 9640 12980
rect 10140 12971 10192 12980
rect 10140 12937 10149 12971
rect 10149 12937 10183 12971
rect 10183 12937 10192 12971
rect 10140 12928 10192 12937
rect 11060 12928 11112 12980
rect 12440 12928 12492 12980
rect 12900 12928 12952 12980
rect 13452 12971 13504 12980
rect 13452 12937 13461 12971
rect 13461 12937 13495 12971
rect 13495 12937 13504 12971
rect 13452 12928 13504 12937
rect 14280 12971 14332 12980
rect 14280 12937 14289 12971
rect 14289 12937 14323 12971
rect 14323 12937 14332 12971
rect 14280 12928 14332 12937
rect 14464 12928 14516 12980
rect 9680 12860 9732 12912
rect 5540 12792 5592 12844
rect 7748 12792 7800 12844
rect 6368 12724 6420 12776
rect 8484 12835 8536 12844
rect 8484 12801 8493 12835
rect 8493 12801 8527 12835
rect 8527 12801 8536 12835
rect 8484 12792 8536 12801
rect 11152 12860 11204 12912
rect 11612 12860 11664 12912
rect 11980 12835 12032 12844
rect 11980 12801 11989 12835
rect 11989 12801 12023 12835
rect 12023 12801 12032 12835
rect 11980 12792 12032 12801
rect 13360 12860 13412 12912
rect 16212 12971 16264 12980
rect 16212 12937 16221 12971
rect 16221 12937 16255 12971
rect 16255 12937 16264 12971
rect 16212 12928 16264 12937
rect 15476 12860 15528 12912
rect 9312 12724 9364 12776
rect 9496 12724 9548 12776
rect 5632 12656 5684 12708
rect 6920 12656 6972 12708
rect 10692 12699 10744 12708
rect 10692 12665 10701 12699
rect 10701 12665 10735 12699
rect 10735 12665 10744 12699
rect 10692 12656 10744 12665
rect 11152 12767 11204 12776
rect 11152 12733 11161 12767
rect 11161 12733 11195 12767
rect 11195 12733 11204 12767
rect 11152 12724 11204 12733
rect 11336 12724 11388 12776
rect 12072 12724 12124 12776
rect 12624 12835 12676 12844
rect 12624 12801 12633 12835
rect 12633 12801 12667 12835
rect 12667 12801 12676 12835
rect 12624 12792 12676 12801
rect 12808 12835 12860 12844
rect 12808 12801 12817 12835
rect 12817 12801 12851 12835
rect 12851 12801 12860 12835
rect 12808 12792 12860 12801
rect 13084 12792 13136 12844
rect 13636 12767 13688 12776
rect 13636 12733 13645 12767
rect 13645 12733 13679 12767
rect 13679 12733 13688 12767
rect 13636 12724 13688 12733
rect 14280 12792 14332 12844
rect 14372 12792 14424 12844
rect 3148 12588 3200 12640
rect 11244 12588 11296 12640
rect 15568 12835 15620 12844
rect 15568 12801 15577 12835
rect 15577 12801 15611 12835
rect 15611 12801 15620 12835
rect 15568 12792 15620 12801
rect 15752 12792 15804 12844
rect 16120 12835 16172 12844
rect 16120 12801 16129 12835
rect 16129 12801 16163 12835
rect 16163 12801 16172 12835
rect 16120 12792 16172 12801
rect 16396 12835 16448 12844
rect 16396 12801 16405 12835
rect 16405 12801 16439 12835
rect 16439 12801 16448 12835
rect 16396 12792 16448 12801
rect 16764 12792 16816 12844
rect 16948 12835 17000 12844
rect 16948 12801 16957 12835
rect 16957 12801 16991 12835
rect 16991 12801 17000 12835
rect 16948 12792 17000 12801
rect 15660 12724 15712 12776
rect 16580 12724 16632 12776
rect 15844 12656 15896 12708
rect 13912 12631 13964 12640
rect 13912 12597 13921 12631
rect 13921 12597 13955 12631
rect 13955 12597 13964 12631
rect 13912 12588 13964 12597
rect 16212 12588 16264 12640
rect 1918 12486 1970 12538
rect 1982 12486 2034 12538
rect 2046 12486 2098 12538
rect 2110 12486 2162 12538
rect 2174 12486 2226 12538
rect 2238 12486 2290 12538
rect 7918 12486 7970 12538
rect 7982 12486 8034 12538
rect 8046 12486 8098 12538
rect 8110 12486 8162 12538
rect 8174 12486 8226 12538
rect 8238 12486 8290 12538
rect 13918 12486 13970 12538
rect 13982 12486 14034 12538
rect 14046 12486 14098 12538
rect 14110 12486 14162 12538
rect 14174 12486 14226 12538
rect 14238 12486 14290 12538
rect 2320 12384 2372 12436
rect 3424 12384 3476 12436
rect 4068 12427 4120 12436
rect 4068 12393 4077 12427
rect 4077 12393 4111 12427
rect 4111 12393 4120 12427
rect 4068 12384 4120 12393
rect 4712 12384 4764 12436
rect 5632 12384 5684 12436
rect 7104 12427 7156 12436
rect 7104 12393 7113 12427
rect 7113 12393 7147 12427
rect 7147 12393 7156 12427
rect 7104 12384 7156 12393
rect 15568 12384 15620 12436
rect 15752 12384 15804 12436
rect 4252 12316 4304 12368
rect 5172 12316 5224 12368
rect 1400 12180 1452 12232
rect 2504 12180 2556 12232
rect 4988 12248 5040 12300
rect 7656 12316 7708 12368
rect 14464 12248 14516 12300
rect 16212 12248 16264 12300
rect 4160 12180 4212 12232
rect 3700 12112 3752 12164
rect 4528 12180 4580 12232
rect 6184 12223 6236 12232
rect 6184 12189 6193 12223
rect 6193 12189 6227 12223
rect 6227 12189 6236 12223
rect 6184 12180 6236 12189
rect 16948 12248 17000 12300
rect 7564 12155 7616 12164
rect 848 12044 900 12096
rect 4344 12044 4396 12096
rect 7564 12121 7573 12155
rect 7573 12121 7607 12155
rect 7607 12121 7616 12155
rect 7564 12112 7616 12121
rect 16764 12180 16816 12232
rect 6644 12044 6696 12096
rect 12532 12044 12584 12096
rect 13176 12044 13228 12096
rect 15660 12044 15712 12096
rect 16120 12044 16172 12096
rect 2658 11942 2710 11994
rect 2722 11942 2774 11994
rect 2786 11942 2838 11994
rect 2850 11942 2902 11994
rect 2914 11942 2966 11994
rect 2978 11942 3030 11994
rect 8658 11942 8710 11994
rect 8722 11942 8774 11994
rect 8786 11942 8838 11994
rect 8850 11942 8902 11994
rect 8914 11942 8966 11994
rect 8978 11942 9030 11994
rect 14658 11942 14710 11994
rect 14722 11942 14774 11994
rect 14786 11942 14838 11994
rect 14850 11942 14902 11994
rect 14914 11942 14966 11994
rect 14978 11942 15030 11994
rect 3608 11883 3660 11892
rect 3608 11849 3617 11883
rect 3617 11849 3651 11883
rect 3651 11849 3660 11883
rect 3608 11840 3660 11849
rect 4344 11840 4396 11892
rect 5448 11840 5500 11892
rect 6184 11840 6236 11892
rect 7564 11840 7616 11892
rect 3424 11704 3476 11756
rect 4160 11747 4212 11756
rect 4160 11713 4169 11747
rect 4169 11713 4203 11747
rect 4203 11713 4212 11747
rect 4160 11704 4212 11713
rect 4252 11636 4304 11688
rect 3700 11568 3752 11620
rect 4528 11747 4580 11756
rect 4528 11713 4537 11747
rect 4537 11713 4571 11747
rect 4571 11713 4580 11747
rect 4528 11704 4580 11713
rect 4804 11704 4856 11756
rect 6920 11747 6972 11756
rect 6920 11713 6929 11747
rect 6929 11713 6963 11747
rect 6963 11713 6972 11747
rect 6920 11704 6972 11713
rect 7012 11704 7064 11756
rect 12716 11840 12768 11892
rect 13084 11840 13136 11892
rect 8392 11747 8444 11756
rect 8392 11713 8401 11747
rect 8401 11713 8435 11747
rect 8435 11713 8444 11747
rect 8392 11704 8444 11713
rect 8484 11747 8536 11756
rect 8484 11713 8493 11747
rect 8493 11713 8527 11747
rect 8527 11713 8536 11747
rect 8484 11704 8536 11713
rect 8852 11704 8904 11756
rect 11612 11772 11664 11824
rect 8392 11568 8444 11620
rect 9772 11704 9824 11756
rect 9312 11568 9364 11620
rect 10508 11704 10560 11756
rect 10784 11704 10836 11756
rect 12532 11704 12584 11756
rect 12716 11747 12768 11756
rect 12716 11713 12725 11747
rect 12725 11713 12759 11747
rect 12759 11713 12768 11747
rect 12716 11704 12768 11713
rect 12900 11704 12952 11756
rect 15292 11772 15344 11824
rect 11612 11568 11664 11620
rect 12624 11679 12676 11688
rect 12624 11645 12633 11679
rect 12633 11645 12667 11679
rect 12667 11645 12676 11679
rect 12624 11636 12676 11645
rect 14556 11704 14608 11756
rect 15844 11840 15896 11892
rect 16948 11840 17000 11892
rect 16580 11772 16632 11824
rect 13176 11636 13228 11688
rect 13452 11636 13504 11688
rect 15108 11679 15160 11688
rect 15108 11645 15117 11679
rect 15117 11645 15151 11679
rect 15151 11645 15160 11679
rect 15108 11636 15160 11645
rect 15660 11747 15712 11756
rect 15660 11713 15669 11747
rect 15669 11713 15703 11747
rect 15703 11713 15712 11747
rect 15660 11704 15712 11713
rect 15752 11747 15804 11756
rect 15752 11713 15761 11747
rect 15761 11713 15795 11747
rect 15795 11713 15804 11747
rect 15752 11704 15804 11713
rect 16028 11704 16080 11756
rect 16212 11704 16264 11756
rect 16764 11704 16816 11756
rect 16948 11704 17000 11756
rect 11704 11500 11756 11552
rect 12992 11500 13044 11552
rect 13636 11500 13688 11552
rect 15660 11500 15712 11552
rect 17040 11500 17092 11552
rect 1918 11398 1970 11450
rect 1982 11398 2034 11450
rect 2046 11398 2098 11450
rect 2110 11398 2162 11450
rect 2174 11398 2226 11450
rect 2238 11398 2290 11450
rect 7918 11398 7970 11450
rect 7982 11398 8034 11450
rect 8046 11398 8098 11450
rect 8110 11398 8162 11450
rect 8174 11398 8226 11450
rect 8238 11398 8290 11450
rect 13918 11398 13970 11450
rect 13982 11398 14034 11450
rect 14046 11398 14098 11450
rect 14110 11398 14162 11450
rect 14174 11398 14226 11450
rect 14238 11398 14290 11450
rect 1400 11339 1452 11348
rect 1400 11305 1409 11339
rect 1409 11305 1443 11339
rect 1443 11305 1452 11339
rect 1400 11296 1452 11305
rect 4804 11339 4856 11348
rect 4804 11305 4813 11339
rect 4813 11305 4847 11339
rect 4847 11305 4856 11339
rect 4804 11296 4856 11305
rect 5448 11339 5500 11348
rect 5448 11305 5457 11339
rect 5457 11305 5491 11339
rect 5491 11305 5500 11339
rect 5448 11296 5500 11305
rect 10784 11339 10836 11348
rect 10784 11305 10793 11339
rect 10793 11305 10827 11339
rect 10827 11305 10836 11339
rect 10784 11296 10836 11305
rect 15660 11339 15712 11348
rect 15660 11305 15669 11339
rect 15669 11305 15703 11339
rect 15703 11305 15712 11339
rect 15660 11296 15712 11305
rect 3148 11203 3200 11212
rect 3148 11169 3157 11203
rect 3157 11169 3191 11203
rect 3191 11169 3200 11203
rect 3148 11160 3200 11169
rect 3700 11160 3752 11212
rect 6920 11228 6972 11280
rect 8484 11203 8536 11212
rect 8484 11169 8493 11203
rect 8493 11169 8527 11203
rect 8527 11169 8536 11203
rect 8484 11160 8536 11169
rect 10508 11203 10560 11212
rect 10508 11169 10517 11203
rect 10517 11169 10551 11203
rect 10551 11169 10560 11203
rect 10508 11160 10560 11169
rect 11704 11160 11756 11212
rect 12716 11160 12768 11212
rect 12992 11203 13044 11212
rect 12992 11169 13001 11203
rect 13001 11169 13035 11203
rect 13035 11169 13044 11203
rect 12992 11160 13044 11169
rect 14372 11160 14424 11212
rect 16120 11228 16172 11280
rect 2504 10956 2556 11008
rect 7012 11135 7064 11144
rect 7012 11101 7021 11135
rect 7021 11101 7055 11135
rect 7055 11101 7064 11135
rect 7012 11092 7064 11101
rect 8392 11135 8444 11144
rect 8392 11101 8401 11135
rect 8401 11101 8435 11135
rect 8435 11101 8444 11135
rect 8392 11092 8444 11101
rect 8852 11092 8904 11144
rect 6920 11024 6972 11076
rect 8484 11024 8536 11076
rect 11612 11092 11664 11144
rect 12440 11092 12492 11144
rect 13268 11092 13320 11144
rect 13452 11092 13504 11144
rect 15384 11160 15436 11212
rect 10692 10956 10744 11008
rect 13360 11024 13412 11076
rect 13728 11024 13780 11076
rect 15292 11135 15344 11144
rect 15292 11101 15301 11135
rect 15301 11101 15335 11135
rect 15335 11101 15344 11135
rect 15292 11092 15344 11101
rect 17040 11160 17092 11212
rect 15752 11092 15804 11144
rect 16764 11092 16816 11144
rect 16120 11067 16172 11076
rect 16120 11033 16129 11067
rect 16129 11033 16163 11067
rect 16163 11033 16172 11067
rect 16120 11024 16172 11033
rect 16304 11067 16356 11076
rect 16304 11033 16313 11067
rect 16313 11033 16347 11067
rect 16347 11033 16356 11067
rect 16304 11024 16356 11033
rect 2658 10854 2710 10906
rect 2722 10854 2774 10906
rect 2786 10854 2838 10906
rect 2850 10854 2902 10906
rect 2914 10854 2966 10906
rect 2978 10854 3030 10906
rect 8658 10854 8710 10906
rect 8722 10854 8774 10906
rect 8786 10854 8838 10906
rect 8850 10854 8902 10906
rect 8914 10854 8966 10906
rect 8978 10854 9030 10906
rect 14658 10854 14710 10906
rect 14722 10854 14774 10906
rect 14786 10854 14838 10906
rect 14850 10854 14902 10906
rect 14914 10854 14966 10906
rect 14978 10854 15030 10906
rect 1308 10752 1360 10804
rect 15108 10752 15160 10804
rect 6644 10684 6696 10736
rect 16580 10684 16632 10736
rect 1400 10616 1452 10668
rect 6368 10659 6420 10668
rect 6368 10625 6377 10659
rect 6377 10625 6411 10659
rect 6411 10625 6420 10659
rect 6368 10616 6420 10625
rect 11612 10616 11664 10668
rect 5724 10548 5776 10600
rect 7104 10548 7156 10600
rect 10784 10548 10836 10600
rect 10968 10548 11020 10600
rect 15752 10616 15804 10668
rect 15200 10548 15252 10600
rect 15660 10548 15712 10600
rect 16672 10659 16724 10668
rect 16672 10625 16681 10659
rect 16681 10625 16715 10659
rect 16715 10625 16724 10659
rect 16672 10616 16724 10625
rect 16764 10659 16816 10668
rect 16764 10625 16773 10659
rect 16773 10625 16807 10659
rect 16807 10625 16816 10659
rect 16764 10616 16816 10625
rect 16948 10591 17000 10600
rect 16948 10557 16957 10591
rect 16957 10557 16991 10591
rect 16991 10557 17000 10591
rect 16948 10548 17000 10557
rect 17040 10480 17092 10532
rect 9680 10412 9732 10464
rect 10876 10412 10928 10464
rect 16948 10412 17000 10464
rect 1918 10310 1970 10362
rect 1982 10310 2034 10362
rect 2046 10310 2098 10362
rect 2110 10310 2162 10362
rect 2174 10310 2226 10362
rect 2238 10310 2290 10362
rect 7918 10310 7970 10362
rect 7982 10310 8034 10362
rect 8046 10310 8098 10362
rect 8110 10310 8162 10362
rect 8174 10310 8226 10362
rect 8238 10310 8290 10362
rect 13918 10310 13970 10362
rect 13982 10310 14034 10362
rect 14046 10310 14098 10362
rect 14110 10310 14162 10362
rect 14174 10310 14226 10362
rect 14238 10310 14290 10362
rect 1400 10251 1452 10260
rect 1400 10217 1409 10251
rect 1409 10217 1443 10251
rect 1443 10217 1452 10251
rect 1400 10208 1452 10217
rect 6644 10251 6696 10260
rect 6644 10217 6653 10251
rect 6653 10217 6687 10251
rect 6687 10217 6696 10251
rect 6644 10208 6696 10217
rect 12716 10208 12768 10260
rect 13268 10208 13320 10260
rect 3884 10183 3936 10192
rect 3884 10149 3893 10183
rect 3893 10149 3927 10183
rect 3927 10149 3936 10183
rect 3884 10140 3936 10149
rect 9772 10140 9824 10192
rect 10784 10140 10836 10192
rect 3148 10047 3200 10056
rect 3148 10013 3157 10047
rect 3157 10013 3191 10047
rect 3191 10013 3200 10047
rect 3148 10004 3200 10013
rect 2412 9936 2464 9988
rect 4252 9979 4304 9988
rect 4252 9945 4261 9979
rect 4261 9945 4295 9979
rect 4295 9945 4304 9979
rect 4252 9936 4304 9945
rect 2504 9868 2556 9920
rect 9772 9936 9824 9988
rect 10048 10047 10100 10056
rect 10048 10013 10057 10047
rect 10057 10013 10091 10047
rect 10091 10013 10100 10047
rect 10048 10004 10100 10013
rect 10692 10115 10744 10124
rect 10692 10081 10701 10115
rect 10701 10081 10735 10115
rect 10735 10081 10744 10115
rect 10692 10072 10744 10081
rect 10876 10047 10928 10056
rect 10876 10013 10885 10047
rect 10885 10013 10919 10047
rect 10919 10013 10928 10047
rect 10876 10004 10928 10013
rect 11612 9936 11664 9988
rect 12900 10140 12952 10192
rect 13636 10140 13688 10192
rect 14096 10140 14148 10192
rect 14464 10140 14516 10192
rect 15200 10208 15252 10260
rect 16856 10208 16908 10260
rect 12532 10047 12584 10056
rect 12532 10013 12541 10047
rect 12541 10013 12575 10047
rect 12575 10013 12584 10047
rect 12532 10004 12584 10013
rect 13452 10072 13504 10124
rect 12716 10004 12768 10056
rect 13084 10047 13136 10056
rect 13084 10013 13093 10047
rect 13093 10013 13127 10047
rect 13127 10013 13136 10047
rect 13084 10004 13136 10013
rect 13544 10004 13596 10056
rect 13912 10004 13964 10056
rect 14556 10047 14608 10056
rect 14556 10013 14565 10047
rect 14565 10013 14599 10047
rect 14599 10013 14608 10047
rect 14556 10004 14608 10013
rect 15752 10072 15804 10124
rect 12992 9936 13044 9988
rect 13452 9936 13504 9988
rect 15292 10004 15344 10056
rect 15568 10004 15620 10056
rect 15660 10004 15712 10056
rect 16580 10140 16632 10192
rect 16672 10183 16724 10192
rect 16672 10149 16681 10183
rect 16681 10149 16715 10183
rect 16715 10149 16724 10183
rect 16672 10140 16724 10149
rect 16948 10047 17000 10056
rect 16948 10013 16957 10047
rect 16957 10013 16991 10047
rect 16991 10013 17000 10047
rect 16948 10004 17000 10013
rect 17040 10047 17092 10056
rect 17040 10013 17049 10047
rect 17049 10013 17083 10047
rect 17083 10013 17092 10047
rect 17040 10004 17092 10013
rect 17132 10004 17184 10056
rect 10048 9868 10100 9920
rect 10968 9868 11020 9920
rect 12532 9868 12584 9920
rect 12716 9911 12768 9920
rect 12716 9877 12725 9911
rect 12725 9877 12759 9911
rect 12759 9877 12768 9911
rect 12716 9868 12768 9877
rect 12900 9911 12952 9920
rect 12900 9877 12909 9911
rect 12909 9877 12943 9911
rect 12943 9877 12952 9911
rect 12900 9868 12952 9877
rect 14556 9868 14608 9920
rect 15568 9868 15620 9920
rect 16580 9911 16632 9920
rect 16580 9877 16589 9911
rect 16589 9877 16623 9911
rect 16623 9877 16632 9911
rect 16580 9868 16632 9877
rect 2658 9766 2710 9818
rect 2722 9766 2774 9818
rect 2786 9766 2838 9818
rect 2850 9766 2902 9818
rect 2914 9766 2966 9818
rect 2978 9766 3030 9818
rect 8658 9766 8710 9818
rect 8722 9766 8774 9818
rect 8786 9766 8838 9818
rect 8850 9766 8902 9818
rect 8914 9766 8966 9818
rect 8978 9766 9030 9818
rect 14658 9766 14710 9818
rect 14722 9766 14774 9818
rect 14786 9766 14838 9818
rect 14850 9766 14902 9818
rect 14914 9766 14966 9818
rect 14978 9766 15030 9818
rect 3884 9664 3936 9716
rect 2412 9639 2464 9648
rect 2412 9605 2421 9639
rect 2421 9605 2455 9639
rect 2455 9605 2464 9639
rect 2412 9596 2464 9605
rect 1400 9528 1452 9580
rect 2504 9571 2556 9580
rect 2504 9537 2513 9571
rect 2513 9537 2547 9571
rect 2547 9537 2556 9571
rect 2504 9528 2556 9537
rect 3424 9571 3476 9580
rect 3424 9537 3433 9571
rect 3433 9537 3467 9571
rect 3467 9537 3476 9571
rect 3424 9528 3476 9537
rect 3516 9571 3568 9580
rect 3516 9537 3525 9571
rect 3525 9537 3559 9571
rect 3559 9537 3568 9571
rect 3516 9528 3568 9537
rect 3976 9528 4028 9580
rect 4068 9571 4120 9580
rect 4068 9537 4077 9571
rect 4077 9537 4111 9571
rect 4111 9537 4120 9571
rect 4068 9528 4120 9537
rect 4712 9571 4764 9580
rect 4712 9537 4721 9571
rect 4721 9537 4755 9571
rect 4755 9537 4764 9571
rect 4712 9528 4764 9537
rect 4896 9571 4948 9580
rect 4896 9537 4905 9571
rect 4905 9537 4939 9571
rect 4939 9537 4948 9571
rect 4896 9528 4948 9537
rect 5080 9528 5132 9580
rect 2412 9460 2464 9512
rect 3700 9460 3752 9512
rect 4160 9503 4212 9512
rect 4160 9469 4169 9503
rect 4169 9469 4203 9503
rect 4203 9469 4212 9503
rect 4160 9460 4212 9469
rect 4436 9460 4488 9512
rect 5724 9596 5776 9648
rect 9680 9596 9732 9648
rect 1308 9392 1360 9444
rect 3148 9392 3200 9444
rect 8392 9460 8444 9512
rect 9772 9571 9824 9580
rect 9772 9537 9781 9571
rect 9781 9537 9815 9571
rect 9815 9537 9824 9571
rect 9772 9528 9824 9537
rect 10048 9460 10100 9512
rect 10692 9528 10744 9580
rect 11336 9528 11388 9580
rect 12624 9664 12676 9716
rect 13084 9664 13136 9716
rect 11980 9503 12032 9512
rect 11980 9469 11989 9503
rect 11989 9469 12023 9503
rect 12023 9469 12032 9503
rect 11980 9460 12032 9469
rect 14188 9596 14240 9648
rect 3424 9324 3476 9376
rect 4160 9324 4212 9376
rect 5264 9367 5316 9376
rect 5264 9333 5273 9367
rect 5273 9333 5307 9367
rect 5307 9333 5316 9367
rect 5264 9324 5316 9333
rect 7288 9324 7340 9376
rect 8668 9324 8720 9376
rect 9220 9324 9272 9376
rect 9496 9324 9548 9376
rect 11888 9367 11940 9376
rect 11888 9333 11897 9367
rect 11897 9333 11931 9367
rect 11931 9333 11940 9367
rect 11888 9324 11940 9333
rect 12072 9367 12124 9376
rect 12072 9333 12081 9367
rect 12081 9333 12115 9367
rect 12115 9333 12124 9367
rect 12072 9324 12124 9333
rect 12532 9571 12584 9580
rect 12532 9537 12541 9571
rect 12541 9537 12575 9571
rect 12575 9537 12584 9571
rect 12532 9528 12584 9537
rect 12624 9571 12676 9580
rect 12624 9537 12633 9571
rect 12633 9537 12667 9571
rect 12667 9537 12676 9571
rect 12624 9528 12676 9537
rect 12900 9571 12952 9580
rect 12900 9537 12909 9571
rect 12909 9537 12943 9571
rect 12943 9537 12952 9571
rect 12900 9528 12952 9537
rect 13084 9571 13136 9580
rect 13084 9537 13093 9571
rect 13093 9537 13127 9571
rect 13127 9537 13136 9571
rect 13084 9528 13136 9537
rect 13452 9571 13504 9580
rect 13452 9537 13461 9571
rect 13461 9537 13495 9571
rect 13495 9537 13504 9571
rect 13452 9528 13504 9537
rect 13820 9528 13872 9580
rect 15476 9664 15528 9716
rect 12992 9460 13044 9512
rect 13176 9503 13228 9512
rect 13176 9469 13185 9503
rect 13185 9469 13219 9503
rect 13219 9469 13228 9503
rect 13176 9460 13228 9469
rect 14924 9528 14976 9580
rect 15200 9596 15252 9648
rect 15384 9577 15436 9586
rect 15384 9543 15389 9577
rect 15389 9543 15423 9577
rect 15423 9543 15436 9577
rect 15384 9534 15436 9543
rect 15476 9528 15528 9580
rect 15568 9571 15620 9580
rect 15568 9537 15577 9571
rect 15577 9537 15611 9571
rect 15611 9537 15620 9571
rect 15568 9528 15620 9537
rect 15660 9571 15712 9580
rect 15660 9537 15669 9571
rect 15669 9537 15703 9571
rect 15703 9537 15712 9571
rect 15660 9528 15712 9537
rect 15752 9571 15804 9580
rect 15752 9537 15761 9571
rect 15761 9537 15795 9571
rect 15795 9537 15804 9571
rect 15752 9528 15804 9537
rect 16120 9596 16172 9648
rect 16580 9528 16632 9580
rect 16856 9571 16908 9580
rect 16856 9537 16865 9571
rect 16865 9537 16899 9571
rect 16899 9537 16908 9571
rect 16856 9528 16908 9537
rect 17224 9571 17276 9580
rect 17224 9537 17233 9571
rect 17233 9537 17267 9571
rect 17267 9537 17276 9571
rect 17224 9528 17276 9537
rect 12808 9392 12860 9444
rect 13360 9392 13412 9444
rect 12440 9324 12492 9376
rect 13452 9324 13504 9376
rect 14004 9324 14056 9376
rect 14464 9503 14516 9512
rect 14464 9469 14473 9503
rect 14473 9469 14507 9503
rect 14507 9469 14516 9503
rect 14464 9460 14516 9469
rect 15108 9460 15160 9512
rect 14924 9392 14976 9444
rect 14556 9324 14608 9376
rect 15016 9324 15068 9376
rect 15292 9503 15344 9512
rect 15292 9469 15301 9503
rect 15301 9469 15335 9503
rect 15335 9469 15344 9503
rect 15292 9460 15344 9469
rect 17132 9460 17184 9512
rect 16120 9324 16172 9376
rect 17040 9324 17092 9376
rect 1918 9222 1970 9274
rect 1982 9222 2034 9274
rect 2046 9222 2098 9274
rect 2110 9222 2162 9274
rect 2174 9222 2226 9274
rect 2238 9222 2290 9274
rect 7918 9222 7970 9274
rect 7982 9222 8034 9274
rect 8046 9222 8098 9274
rect 8110 9222 8162 9274
rect 8174 9222 8226 9274
rect 8238 9222 8290 9274
rect 13918 9222 13970 9274
rect 13982 9222 14034 9274
rect 14046 9222 14098 9274
rect 14110 9222 14162 9274
rect 14174 9222 14226 9274
rect 14238 9222 14290 9274
rect 1400 9163 1452 9172
rect 1400 9129 1409 9163
rect 1409 9129 1443 9163
rect 1443 9129 1452 9163
rect 1400 9120 1452 9129
rect 3516 9120 3568 9172
rect 4160 9120 4212 9172
rect 4252 9120 4304 9172
rect 6920 9120 6972 9172
rect 8392 9120 8444 9172
rect 8484 9120 8536 9172
rect 3148 9027 3200 9036
rect 3148 8993 3157 9027
rect 3157 8993 3191 9027
rect 3191 8993 3200 9027
rect 3148 8984 3200 8993
rect 3976 8916 4028 8968
rect 12072 9120 12124 9172
rect 12624 9163 12676 9172
rect 12624 9129 12633 9163
rect 12633 9129 12667 9163
rect 12667 9129 12676 9163
rect 12624 9120 12676 9129
rect 14556 9120 14608 9172
rect 14924 9120 14976 9172
rect 4712 8984 4764 9036
rect 4896 8916 4948 8968
rect 2228 8848 2280 8900
rect 4068 8891 4120 8900
rect 4068 8857 4077 8891
rect 4077 8857 4111 8891
rect 4111 8857 4120 8891
rect 4068 8848 4120 8857
rect 5264 8848 5316 8900
rect 5540 8959 5592 8968
rect 5540 8925 5549 8959
rect 5549 8925 5583 8959
rect 5583 8925 5592 8959
rect 5540 8916 5592 8925
rect 5632 8916 5684 8968
rect 9680 9052 9732 9104
rect 13360 9052 13412 9104
rect 5724 8848 5776 8900
rect 7288 8959 7340 8968
rect 7288 8925 7297 8959
rect 7297 8925 7331 8959
rect 7331 8925 7340 8959
rect 7288 8916 7340 8925
rect 9220 8984 9272 9036
rect 11980 8984 12032 9036
rect 7380 8848 7432 8900
rect 8668 8959 8720 8968
rect 8668 8925 8677 8959
rect 8677 8925 8711 8959
rect 8711 8925 8720 8959
rect 8668 8916 8720 8925
rect 12808 8984 12860 9036
rect 12716 8916 12768 8968
rect 13176 8916 13228 8968
rect 15200 9052 15252 9104
rect 15292 9052 15344 9104
rect 14464 8984 14516 9036
rect 17224 9052 17276 9104
rect 17040 9027 17092 9036
rect 17040 8993 17049 9027
rect 17049 8993 17083 9027
rect 17083 8993 17092 9027
rect 17040 8984 17092 8993
rect 15016 8959 15068 8968
rect 15016 8925 15025 8959
rect 15025 8925 15059 8959
rect 15059 8925 15068 8959
rect 15016 8916 15068 8925
rect 15108 8959 15160 8968
rect 15108 8925 15117 8959
rect 15117 8925 15151 8959
rect 15151 8925 15160 8959
rect 15108 8916 15160 8925
rect 15200 8916 15252 8968
rect 15844 8916 15896 8968
rect 9496 8848 9548 8900
rect 14556 8848 14608 8900
rect 16856 8916 16908 8968
rect 17132 8959 17184 8968
rect 17132 8925 17141 8959
rect 17141 8925 17175 8959
rect 17175 8925 17184 8959
rect 17132 8916 17184 8925
rect 16764 8848 16816 8900
rect 3056 8780 3108 8832
rect 3976 8823 4028 8832
rect 3976 8789 3985 8823
rect 3985 8789 4019 8823
rect 4019 8789 4028 8823
rect 3976 8780 4028 8789
rect 12716 8780 12768 8832
rect 13268 8780 13320 8832
rect 15108 8780 15160 8832
rect 16396 8823 16448 8832
rect 16396 8789 16405 8823
rect 16405 8789 16439 8823
rect 16439 8789 16448 8823
rect 16396 8780 16448 8789
rect 2658 8678 2710 8730
rect 2722 8678 2774 8730
rect 2786 8678 2838 8730
rect 2850 8678 2902 8730
rect 2914 8678 2966 8730
rect 2978 8678 3030 8730
rect 8658 8678 8710 8730
rect 8722 8678 8774 8730
rect 8786 8678 8838 8730
rect 8850 8678 8902 8730
rect 8914 8678 8966 8730
rect 8978 8678 9030 8730
rect 14658 8678 14710 8730
rect 14722 8678 14774 8730
rect 14786 8678 14838 8730
rect 14850 8678 14902 8730
rect 14914 8678 14966 8730
rect 14978 8678 15030 8730
rect 1308 8576 1360 8628
rect 2228 8619 2280 8628
rect 2228 8585 2237 8619
rect 2237 8585 2271 8619
rect 2271 8585 2280 8619
rect 2228 8576 2280 8585
rect 5264 8576 5316 8628
rect 5724 8619 5776 8628
rect 5724 8585 5733 8619
rect 5733 8585 5767 8619
rect 5767 8585 5776 8619
rect 5724 8576 5776 8585
rect 9220 8619 9272 8628
rect 9220 8585 9229 8619
rect 9229 8585 9263 8619
rect 9263 8585 9272 8619
rect 9220 8576 9272 8585
rect 11520 8576 11572 8628
rect 1584 8483 1636 8492
rect 1584 8449 1593 8483
rect 1593 8449 1627 8483
rect 1627 8449 1636 8483
rect 1584 8440 1636 8449
rect 2412 8440 2464 8492
rect 4160 8440 4212 8492
rect 5172 8483 5224 8492
rect 5172 8449 5200 8483
rect 5200 8449 5224 8483
rect 5172 8440 5224 8449
rect 5356 8483 5408 8492
rect 5356 8449 5365 8483
rect 5365 8449 5399 8483
rect 5399 8449 5408 8483
rect 5356 8440 5408 8449
rect 5632 8483 5684 8492
rect 5632 8449 5641 8483
rect 5641 8449 5675 8483
rect 5675 8449 5684 8483
rect 5632 8440 5684 8449
rect 3056 8372 3108 8424
rect 3424 8372 3476 8424
rect 3976 8372 4028 8424
rect 5172 8236 5224 8288
rect 7196 8483 7248 8492
rect 7196 8449 7205 8483
rect 7205 8449 7239 8483
rect 7239 8449 7248 8483
rect 7196 8440 7248 8449
rect 7472 8483 7524 8492
rect 7472 8449 7481 8483
rect 7481 8449 7515 8483
rect 7515 8449 7524 8483
rect 7472 8440 7524 8449
rect 7656 8483 7708 8492
rect 7656 8449 7665 8483
rect 7665 8449 7699 8483
rect 7699 8449 7708 8483
rect 7656 8440 7708 8449
rect 11888 8508 11940 8560
rect 12256 8508 12308 8560
rect 9588 8483 9640 8492
rect 9588 8449 9597 8483
rect 9597 8449 9631 8483
rect 9631 8449 9640 8483
rect 9588 8440 9640 8449
rect 9680 8483 9732 8492
rect 9680 8449 9689 8483
rect 9689 8449 9723 8483
rect 9723 8449 9732 8483
rect 9680 8440 9732 8449
rect 11336 8440 11388 8492
rect 17132 8576 17184 8628
rect 13084 8440 13136 8492
rect 9956 8372 10008 8424
rect 12072 8415 12124 8424
rect 12072 8381 12081 8415
rect 12081 8381 12115 8415
rect 12115 8381 12124 8415
rect 12072 8372 12124 8381
rect 7380 8304 7432 8356
rect 11612 8347 11664 8356
rect 11612 8313 11621 8347
rect 11621 8313 11655 8347
rect 11655 8313 11664 8347
rect 11612 8304 11664 8313
rect 10140 8236 10192 8288
rect 12440 8279 12492 8288
rect 12440 8245 12449 8279
rect 12449 8245 12483 8279
rect 12483 8245 12492 8279
rect 12440 8236 12492 8245
rect 1918 8134 1970 8186
rect 1982 8134 2034 8186
rect 2046 8134 2098 8186
rect 2110 8134 2162 8186
rect 2174 8134 2226 8186
rect 2238 8134 2290 8186
rect 7918 8134 7970 8186
rect 7982 8134 8034 8186
rect 8046 8134 8098 8186
rect 8110 8134 8162 8186
rect 8174 8134 8226 8186
rect 8238 8134 8290 8186
rect 13918 8134 13970 8186
rect 13982 8134 14034 8186
rect 14046 8134 14098 8186
rect 14110 8134 14162 8186
rect 14174 8134 14226 8186
rect 14238 8134 14290 8186
rect 1584 8032 1636 8084
rect 7472 8032 7524 8084
rect 5540 8007 5592 8016
rect 5540 7973 5549 8007
rect 5549 7973 5583 8007
rect 5583 7973 5592 8007
rect 5540 7964 5592 7973
rect 7196 8007 7248 8016
rect 7196 7973 7205 8007
rect 7205 7973 7239 8007
rect 7239 7973 7248 8007
rect 7196 7964 7248 7973
rect 7380 8007 7432 8016
rect 7380 7973 7389 8007
rect 7389 7973 7423 8007
rect 7423 7973 7432 8007
rect 7380 7964 7432 7973
rect 7656 7964 7708 8016
rect 3148 7939 3200 7948
rect 3148 7905 3157 7939
rect 3157 7905 3191 7939
rect 3191 7905 3200 7939
rect 3148 7896 3200 7905
rect 5356 7896 5408 7948
rect 9956 8075 10008 8084
rect 9956 8041 9965 8075
rect 9965 8041 9999 8075
rect 9999 8041 10008 8075
rect 9956 8032 10008 8041
rect 10140 8032 10192 8084
rect 9680 7964 9732 8016
rect 5172 7871 5224 7880
rect 5172 7837 5181 7871
rect 5181 7837 5215 7871
rect 5215 7837 5224 7871
rect 5172 7828 5224 7837
rect 7380 7828 7432 7880
rect 2320 7760 2372 7812
rect 3424 7760 3476 7812
rect 7840 7828 7892 7880
rect 9956 7896 10008 7948
rect 11060 7939 11112 7948
rect 11060 7905 11069 7939
rect 11069 7905 11103 7939
rect 11103 7905 11112 7939
rect 11060 7896 11112 7905
rect 11796 7896 11848 7948
rect 12072 7896 12124 7948
rect 9496 7828 9548 7880
rect 12440 7828 12492 7880
rect 14464 7828 14516 7880
rect 15752 7871 15804 7880
rect 15752 7837 15761 7871
rect 15761 7837 15795 7871
rect 15795 7837 15804 7871
rect 15752 7828 15804 7837
rect 15936 7871 15988 7880
rect 15936 7837 15949 7871
rect 15949 7837 15988 7871
rect 15936 7828 15988 7837
rect 10140 7760 10192 7812
rect 14372 7760 14424 7812
rect 14556 7692 14608 7744
rect 16212 7692 16264 7744
rect 16488 7692 16540 7744
rect 2658 7590 2710 7642
rect 2722 7590 2774 7642
rect 2786 7590 2838 7642
rect 2850 7590 2902 7642
rect 2914 7590 2966 7642
rect 2978 7590 3030 7642
rect 8658 7590 8710 7642
rect 8722 7590 8774 7642
rect 8786 7590 8838 7642
rect 8850 7590 8902 7642
rect 8914 7590 8966 7642
rect 8978 7590 9030 7642
rect 14658 7590 14710 7642
rect 14722 7590 14774 7642
rect 14786 7590 14838 7642
rect 14850 7590 14902 7642
rect 14914 7590 14966 7642
rect 14978 7590 15030 7642
rect 1308 7488 1360 7540
rect 2320 7531 2372 7540
rect 2320 7497 2329 7531
rect 2329 7497 2363 7531
rect 2363 7497 2372 7531
rect 2320 7488 2372 7497
rect 9496 7531 9548 7540
rect 9496 7497 9505 7531
rect 9505 7497 9539 7531
rect 9539 7497 9548 7531
rect 9496 7488 9548 7497
rect 9588 7531 9640 7540
rect 9588 7497 9597 7531
rect 9597 7497 9631 7531
rect 9631 7497 9640 7531
rect 9588 7488 9640 7497
rect 10140 7531 10192 7540
rect 10140 7497 10149 7531
rect 10149 7497 10183 7531
rect 10183 7497 10192 7531
rect 10140 7488 10192 7497
rect 15752 7488 15804 7540
rect 1584 7395 1636 7404
rect 1584 7361 1593 7395
rect 1593 7361 1627 7395
rect 1627 7361 1636 7395
rect 1584 7352 1636 7361
rect 2412 7395 2464 7404
rect 2412 7361 2421 7395
rect 2421 7361 2455 7395
rect 2455 7361 2464 7395
rect 2412 7352 2464 7361
rect 3884 7352 3936 7404
rect 3424 7327 3476 7336
rect 3424 7293 3433 7327
rect 3433 7293 3467 7327
rect 3467 7293 3476 7327
rect 3424 7284 3476 7293
rect 4804 7352 4856 7404
rect 5816 7352 5868 7404
rect 12440 7463 12492 7472
rect 12440 7429 12449 7463
rect 12449 7429 12483 7463
rect 12483 7429 12492 7463
rect 12440 7420 12492 7429
rect 15108 7420 15160 7472
rect 9772 7395 9824 7404
rect 9772 7361 9781 7395
rect 9781 7361 9815 7395
rect 9815 7361 9824 7395
rect 9772 7352 9824 7361
rect 9956 7395 10008 7404
rect 9956 7361 9965 7395
rect 9965 7361 9999 7395
rect 9999 7361 10008 7395
rect 9956 7352 10008 7361
rect 3792 7216 3844 7268
rect 9864 7216 9916 7268
rect 11060 7352 11112 7404
rect 12164 7395 12216 7404
rect 12164 7361 12173 7395
rect 12173 7361 12207 7395
rect 12207 7361 12216 7395
rect 12164 7352 12216 7361
rect 13544 7352 13596 7404
rect 14372 7352 14424 7404
rect 11244 7284 11296 7336
rect 12072 7284 12124 7336
rect 13636 7284 13688 7336
rect 14464 7284 14516 7336
rect 14648 7327 14700 7336
rect 14648 7293 14657 7327
rect 14657 7293 14691 7327
rect 14691 7293 14700 7327
rect 14648 7284 14700 7293
rect 16488 7352 16540 7404
rect 4712 7191 4764 7200
rect 4712 7157 4721 7191
rect 4721 7157 4755 7191
rect 4755 7157 4764 7191
rect 4712 7148 4764 7157
rect 11428 7216 11480 7268
rect 11520 7148 11572 7200
rect 17224 7191 17276 7200
rect 17224 7157 17233 7191
rect 17233 7157 17267 7191
rect 17267 7157 17276 7191
rect 17224 7148 17276 7157
rect 1918 7046 1970 7098
rect 1982 7046 2034 7098
rect 2046 7046 2098 7098
rect 2110 7046 2162 7098
rect 2174 7046 2226 7098
rect 2238 7046 2290 7098
rect 7918 7046 7970 7098
rect 7982 7046 8034 7098
rect 8046 7046 8098 7098
rect 8110 7046 8162 7098
rect 8174 7046 8226 7098
rect 8238 7046 8290 7098
rect 13918 7046 13970 7098
rect 13982 7046 14034 7098
rect 14046 7046 14098 7098
rect 14110 7046 14162 7098
rect 14174 7046 14226 7098
rect 14238 7046 14290 7098
rect 1584 6944 1636 6996
rect 9956 6944 10008 6996
rect 10600 6944 10652 6996
rect 11060 6987 11112 6996
rect 11060 6953 11069 6987
rect 11069 6953 11103 6987
rect 11103 6953 11112 6987
rect 11060 6944 11112 6953
rect 14372 6944 14424 6996
rect 15200 6944 15252 6996
rect 4804 6876 4856 6928
rect 3148 6851 3200 6860
rect 3148 6817 3157 6851
rect 3157 6817 3191 6851
rect 3191 6817 3200 6851
rect 3148 6808 3200 6817
rect 4160 6808 4212 6860
rect 3792 6783 3844 6792
rect 3792 6749 3801 6783
rect 3801 6749 3835 6783
rect 3835 6749 3844 6783
rect 3792 6740 3844 6749
rect 3884 6783 3936 6792
rect 3884 6749 3893 6783
rect 3893 6749 3927 6783
rect 3927 6749 3936 6783
rect 3884 6740 3936 6749
rect 4712 6740 4764 6792
rect 9128 6808 9180 6860
rect 9772 6808 9824 6860
rect 11428 6808 11480 6860
rect 7472 6740 7524 6792
rect 2320 6672 2372 6724
rect 3608 6672 3660 6724
rect 7564 6715 7616 6724
rect 7564 6681 7573 6715
rect 7573 6681 7607 6715
rect 7607 6681 7616 6715
rect 7564 6672 7616 6681
rect 8576 6604 8628 6656
rect 9404 6783 9456 6792
rect 9404 6749 9413 6783
rect 9413 6749 9447 6783
rect 9447 6749 9456 6783
rect 9404 6740 9456 6749
rect 9312 6672 9364 6724
rect 11520 6783 11572 6792
rect 11520 6749 11529 6783
rect 11529 6749 11563 6783
rect 11563 6749 11572 6783
rect 11520 6740 11572 6749
rect 12256 6808 12308 6860
rect 12624 6808 12676 6860
rect 13544 6808 13596 6860
rect 12072 6783 12124 6792
rect 12072 6749 12081 6783
rect 12081 6749 12115 6783
rect 12115 6749 12124 6783
rect 12072 6740 12124 6749
rect 12164 6740 12216 6792
rect 11612 6672 11664 6724
rect 13084 6740 13136 6792
rect 14372 6851 14424 6860
rect 14372 6817 14381 6851
rect 14381 6817 14415 6851
rect 14415 6817 14424 6851
rect 14372 6808 14424 6817
rect 17224 6851 17276 6860
rect 17224 6817 17233 6851
rect 17233 6817 17267 6851
rect 17267 6817 17276 6851
rect 17224 6808 17276 6817
rect 13820 6783 13872 6792
rect 13820 6749 13829 6783
rect 13829 6749 13863 6783
rect 13863 6749 13872 6783
rect 13820 6740 13872 6749
rect 14004 6740 14056 6792
rect 14556 6783 14608 6792
rect 14556 6749 14565 6783
rect 14565 6749 14599 6783
rect 14599 6749 14608 6783
rect 14556 6740 14608 6749
rect 14740 6783 14792 6792
rect 14740 6749 14749 6783
rect 14749 6749 14783 6783
rect 14783 6749 14792 6783
rect 14740 6740 14792 6749
rect 15016 6740 15068 6792
rect 14648 6672 14700 6724
rect 15200 6783 15252 6792
rect 15200 6749 15209 6783
rect 15209 6749 15243 6783
rect 15243 6749 15252 6783
rect 15200 6740 15252 6749
rect 16212 6740 16264 6792
rect 13912 6604 13964 6656
rect 14372 6604 14424 6656
rect 14740 6604 14792 6656
rect 15108 6604 15160 6656
rect 2658 6502 2710 6554
rect 2722 6502 2774 6554
rect 2786 6502 2838 6554
rect 2850 6502 2902 6554
rect 2914 6502 2966 6554
rect 2978 6502 3030 6554
rect 8658 6502 8710 6554
rect 8722 6502 8774 6554
rect 8786 6502 8838 6554
rect 8850 6502 8902 6554
rect 8914 6502 8966 6554
rect 8978 6502 9030 6554
rect 14658 6502 14710 6554
rect 14722 6502 14774 6554
rect 14786 6502 14838 6554
rect 14850 6502 14902 6554
rect 14914 6502 14966 6554
rect 14978 6502 15030 6554
rect 1308 6400 1360 6452
rect 2320 6443 2372 6452
rect 2320 6409 2329 6443
rect 2329 6409 2363 6443
rect 2363 6409 2372 6443
rect 2320 6400 2372 6409
rect 3792 6400 3844 6452
rect 5816 6443 5868 6452
rect 5816 6409 5825 6443
rect 5825 6409 5859 6443
rect 5859 6409 5868 6443
rect 5816 6400 5868 6409
rect 1584 6307 1636 6316
rect 1584 6273 1593 6307
rect 1593 6273 1627 6307
rect 1627 6273 1636 6307
rect 1584 6264 1636 6273
rect 2412 6307 2464 6316
rect 2412 6273 2421 6307
rect 2421 6273 2455 6307
rect 2455 6273 2464 6307
rect 2412 6264 2464 6273
rect 7656 6332 7708 6384
rect 10140 6400 10192 6452
rect 16304 6400 16356 6452
rect 11888 6332 11940 6384
rect 12256 6332 12308 6384
rect 14280 6332 14332 6384
rect 14372 6332 14424 6384
rect 4252 6307 4304 6316
rect 3608 6239 3660 6248
rect 3608 6205 3617 6239
rect 3617 6205 3651 6239
rect 3651 6205 3660 6239
rect 3608 6196 3660 6205
rect 4252 6273 4261 6307
rect 4261 6273 4295 6307
rect 4295 6273 4304 6307
rect 4252 6264 4304 6273
rect 4344 6307 4396 6316
rect 4344 6273 4353 6307
rect 4353 6273 4387 6307
rect 4387 6273 4396 6307
rect 4344 6264 4396 6273
rect 5908 6264 5960 6316
rect 6736 6307 6788 6316
rect 6736 6273 6745 6307
rect 6745 6273 6779 6307
rect 6779 6273 6788 6307
rect 6736 6264 6788 6273
rect 7380 6264 7432 6316
rect 7748 6196 7800 6248
rect 8392 6264 8444 6316
rect 9864 6307 9916 6316
rect 9864 6273 9873 6307
rect 9873 6273 9907 6307
rect 9907 6273 9916 6307
rect 9864 6264 9916 6273
rect 11612 6264 11664 6316
rect 12624 6307 12676 6316
rect 12624 6273 12636 6307
rect 12636 6273 12670 6307
rect 12670 6273 12676 6307
rect 12624 6264 12676 6273
rect 8576 6239 8628 6248
rect 8576 6205 8585 6239
rect 8585 6205 8619 6239
rect 8619 6205 8628 6239
rect 8576 6196 8628 6205
rect 10140 6239 10192 6248
rect 10140 6205 10149 6239
rect 10149 6205 10183 6239
rect 10183 6205 10192 6239
rect 10140 6196 10192 6205
rect 11796 6239 11848 6248
rect 11796 6205 11805 6239
rect 11805 6205 11839 6239
rect 11839 6205 11848 6239
rect 11796 6196 11848 6205
rect 11520 6128 11572 6180
rect 12440 6196 12492 6248
rect 14556 6264 14608 6316
rect 14832 6264 14884 6316
rect 15936 6128 15988 6180
rect 6368 6060 6420 6112
rect 7840 6060 7892 6112
rect 9956 6103 10008 6112
rect 9956 6069 9965 6103
rect 9965 6069 9999 6103
rect 9999 6069 10008 6103
rect 9956 6060 10008 6069
rect 10048 6103 10100 6112
rect 10048 6069 10057 6103
rect 10057 6069 10091 6103
rect 10091 6069 10100 6103
rect 10048 6060 10100 6069
rect 11888 6060 11940 6112
rect 12624 6060 12676 6112
rect 12808 6060 12860 6112
rect 14372 6060 14424 6112
rect 1918 5958 1970 6010
rect 1982 5958 2034 6010
rect 2046 5958 2098 6010
rect 2110 5958 2162 6010
rect 2174 5958 2226 6010
rect 2238 5958 2290 6010
rect 7918 5958 7970 6010
rect 7982 5958 8034 6010
rect 8046 5958 8098 6010
rect 8110 5958 8162 6010
rect 8174 5958 8226 6010
rect 8238 5958 8290 6010
rect 13918 5958 13970 6010
rect 13982 5958 14034 6010
rect 14046 5958 14098 6010
rect 14110 5958 14162 6010
rect 14174 5958 14226 6010
rect 14238 5958 14290 6010
rect 4252 5899 4304 5908
rect 4252 5865 4261 5899
rect 4261 5865 4295 5899
rect 4295 5865 4304 5899
rect 4252 5856 4304 5865
rect 4344 5856 4396 5908
rect 5908 5856 5960 5908
rect 7656 5899 7708 5908
rect 7656 5865 7665 5899
rect 7665 5865 7699 5899
rect 7699 5865 7708 5899
rect 7656 5856 7708 5865
rect 7748 5856 7800 5908
rect 9956 5856 10008 5908
rect 10416 5856 10468 5908
rect 6368 5831 6420 5840
rect 6368 5797 6377 5831
rect 6377 5797 6411 5831
rect 6411 5797 6420 5831
rect 6368 5788 6420 5797
rect 7104 5788 7156 5840
rect 8208 5788 8260 5840
rect 9220 5788 9272 5840
rect 9864 5788 9916 5840
rect 10232 5788 10284 5840
rect 11152 5899 11204 5908
rect 11152 5865 11161 5899
rect 11161 5865 11195 5899
rect 11195 5865 11204 5899
rect 11152 5856 11204 5865
rect 7380 5720 7432 5772
rect 10600 5788 10652 5840
rect 12624 5856 12676 5908
rect 16212 5899 16264 5908
rect 16212 5865 16221 5899
rect 16221 5865 16255 5899
rect 16255 5865 16264 5899
rect 16212 5856 16264 5865
rect 16488 5899 16540 5908
rect 16488 5865 16497 5899
rect 16497 5865 16531 5899
rect 16531 5865 16540 5899
rect 16488 5856 16540 5865
rect 1492 5652 1544 5704
rect 4436 5695 4488 5704
rect 4436 5661 4445 5695
rect 4445 5661 4479 5695
rect 4479 5661 4488 5695
rect 4436 5652 4488 5661
rect 4620 5652 4672 5704
rect 7472 5695 7524 5704
rect 7472 5661 7481 5695
rect 7481 5661 7515 5695
rect 7515 5661 7524 5695
rect 7472 5652 7524 5661
rect 6644 5627 6696 5636
rect 6644 5593 6653 5627
rect 6653 5593 6687 5627
rect 6687 5593 6696 5627
rect 6644 5584 6696 5593
rect 7932 5695 7984 5704
rect 7932 5661 7941 5695
rect 7941 5661 7975 5695
rect 7975 5661 7984 5695
rect 7932 5652 7984 5661
rect 8116 5695 8168 5704
rect 8116 5661 8125 5695
rect 8125 5661 8159 5695
rect 8159 5661 8168 5695
rect 8116 5652 8168 5661
rect 8208 5695 8260 5704
rect 8208 5661 8217 5695
rect 8217 5661 8251 5695
rect 8251 5661 8260 5695
rect 8208 5652 8260 5661
rect 8300 5695 8352 5704
rect 8300 5661 8309 5695
rect 8309 5661 8343 5695
rect 8343 5661 8352 5695
rect 8300 5652 8352 5661
rect 10324 5720 10376 5772
rect 12164 5788 12216 5840
rect 11888 5720 11940 5772
rect 9128 5584 9180 5636
rect 1400 5559 1452 5568
rect 1400 5525 1409 5559
rect 1409 5525 1443 5559
rect 1443 5525 1452 5559
rect 1400 5516 1452 5525
rect 4160 5516 4212 5568
rect 7196 5516 7248 5568
rect 7564 5516 7616 5568
rect 8116 5516 8168 5568
rect 8484 5516 8536 5568
rect 9772 5695 9824 5704
rect 9772 5661 9781 5695
rect 9781 5661 9815 5695
rect 9815 5661 9824 5695
rect 9772 5652 9824 5661
rect 11796 5652 11848 5704
rect 9772 5516 9824 5568
rect 10324 5516 10376 5568
rect 10692 5627 10744 5636
rect 10692 5593 10701 5627
rect 10701 5593 10735 5627
rect 10735 5593 10744 5627
rect 10692 5584 10744 5593
rect 12256 5584 12308 5636
rect 12348 5627 12400 5636
rect 12348 5593 12357 5627
rect 12357 5593 12391 5627
rect 12391 5593 12400 5627
rect 12348 5584 12400 5593
rect 12624 5695 12676 5704
rect 12624 5661 12633 5695
rect 12633 5661 12667 5695
rect 12667 5661 12676 5695
rect 12624 5652 12676 5661
rect 12900 5763 12952 5772
rect 12900 5729 12909 5763
rect 12909 5729 12943 5763
rect 12943 5729 12952 5763
rect 12900 5720 12952 5729
rect 13452 5720 13504 5772
rect 14280 5788 14332 5840
rect 13728 5763 13780 5772
rect 13728 5729 13737 5763
rect 13737 5729 13771 5763
rect 13771 5729 13780 5763
rect 13728 5720 13780 5729
rect 14648 5720 14700 5772
rect 14832 5720 14884 5772
rect 15568 5763 15620 5772
rect 15568 5729 15577 5763
rect 15577 5729 15611 5763
rect 15611 5729 15620 5763
rect 15568 5720 15620 5729
rect 15384 5695 15436 5704
rect 15384 5661 15393 5695
rect 15393 5661 15427 5695
rect 15427 5661 15436 5695
rect 15384 5652 15436 5661
rect 16580 5788 16632 5840
rect 16396 5720 16448 5772
rect 16672 5763 16724 5772
rect 16672 5729 16681 5763
rect 16681 5729 16715 5763
rect 16715 5729 16724 5763
rect 16672 5720 16724 5729
rect 13452 5627 13504 5636
rect 13452 5593 13461 5627
rect 13461 5593 13495 5627
rect 13495 5593 13504 5627
rect 13452 5584 13504 5593
rect 16304 5627 16356 5636
rect 16304 5593 16313 5627
rect 16313 5593 16347 5627
rect 16347 5593 16356 5627
rect 16304 5584 16356 5593
rect 10876 5516 10928 5568
rect 11060 5516 11112 5568
rect 14096 5559 14148 5568
rect 14096 5525 14105 5559
rect 14105 5525 14139 5559
rect 14139 5525 14148 5559
rect 14096 5516 14148 5525
rect 2658 5414 2710 5466
rect 2722 5414 2774 5466
rect 2786 5414 2838 5466
rect 2850 5414 2902 5466
rect 2914 5414 2966 5466
rect 2978 5414 3030 5466
rect 8658 5414 8710 5466
rect 8722 5414 8774 5466
rect 8786 5414 8838 5466
rect 8850 5414 8902 5466
rect 8914 5414 8966 5466
rect 8978 5414 9030 5466
rect 14658 5414 14710 5466
rect 14722 5414 14774 5466
rect 14786 5414 14838 5466
rect 14850 5414 14902 5466
rect 14914 5414 14966 5466
rect 14978 5414 15030 5466
rect 1584 5312 1636 5364
rect 5816 5312 5868 5364
rect 2320 5244 2372 5296
rect 4436 5244 4488 5296
rect 3148 5219 3200 5228
rect 3148 5185 3157 5219
rect 3157 5185 3191 5219
rect 3191 5185 3200 5219
rect 3148 5176 3200 5185
rect 4160 5176 4212 5228
rect 4620 5219 4672 5228
rect 4620 5185 4628 5219
rect 4628 5185 4662 5219
rect 4662 5185 4672 5219
rect 4620 5176 4672 5185
rect 5908 5287 5960 5296
rect 5908 5253 5917 5287
rect 5917 5253 5951 5287
rect 5951 5253 5960 5287
rect 5908 5244 5960 5253
rect 8300 5312 8352 5364
rect 8668 5312 8720 5364
rect 9220 5312 9272 5364
rect 10324 5312 10376 5364
rect 11704 5312 11756 5364
rect 5448 5219 5500 5228
rect 5448 5185 5457 5219
rect 5457 5185 5491 5219
rect 5491 5185 5500 5219
rect 5448 5176 5500 5185
rect 7196 5219 7248 5228
rect 7196 5185 7205 5219
rect 7205 5185 7239 5219
rect 7239 5185 7248 5219
rect 7196 5176 7248 5185
rect 7472 5176 7524 5228
rect 11152 5244 11204 5296
rect 9128 5176 9180 5228
rect 10140 5176 10192 5228
rect 10416 5219 10468 5228
rect 10416 5185 10425 5219
rect 10425 5185 10459 5219
rect 10459 5185 10468 5219
rect 10416 5176 10468 5185
rect 10508 5176 10560 5228
rect 10692 5219 10744 5228
rect 10692 5185 10701 5219
rect 10701 5185 10735 5219
rect 10735 5185 10744 5219
rect 10692 5176 10744 5185
rect 10784 5219 10836 5228
rect 10784 5185 10793 5219
rect 10793 5185 10827 5219
rect 10827 5185 10836 5219
rect 10784 5176 10836 5185
rect 13728 5312 13780 5364
rect 13820 5312 13872 5364
rect 14096 5244 14148 5296
rect 5908 5108 5960 5160
rect 7380 5151 7432 5160
rect 7380 5117 7389 5151
rect 7389 5117 7423 5151
rect 7423 5117 7432 5151
rect 7380 5108 7432 5117
rect 7656 5108 7708 5160
rect 9220 5108 9272 5160
rect 9496 5108 9548 5160
rect 12808 5219 12860 5228
rect 12808 5185 12817 5219
rect 12817 5185 12851 5219
rect 12851 5185 12860 5219
rect 12808 5176 12860 5185
rect 12532 5108 12584 5160
rect 14280 5219 14332 5228
rect 14280 5185 14289 5219
rect 14289 5185 14323 5219
rect 14323 5185 14332 5219
rect 14280 5176 14332 5185
rect 14372 5219 14424 5228
rect 14372 5185 14381 5219
rect 14381 5185 14415 5219
rect 14415 5185 14424 5219
rect 14372 5176 14424 5185
rect 14556 5176 14608 5228
rect 15292 5219 15344 5228
rect 13728 5108 13780 5160
rect 15292 5185 15323 5219
rect 15323 5185 15344 5219
rect 15292 5176 15344 5185
rect 16304 5312 16356 5364
rect 15936 5244 15988 5296
rect 16028 5219 16080 5228
rect 16028 5185 16037 5219
rect 16037 5185 16071 5219
rect 16071 5185 16080 5219
rect 16028 5176 16080 5185
rect 7196 5083 7248 5092
rect 7196 5049 7205 5083
rect 7205 5049 7239 5083
rect 7239 5049 7248 5083
rect 7196 5040 7248 5049
rect 5816 4972 5868 5024
rect 6644 4972 6696 5024
rect 10968 5040 11020 5092
rect 8668 5015 8720 5024
rect 8668 4981 8677 5015
rect 8677 4981 8711 5015
rect 8711 4981 8720 5015
rect 8668 4972 8720 4981
rect 9312 4972 9364 5024
rect 10232 5015 10284 5024
rect 10232 4981 10241 5015
rect 10241 4981 10275 5015
rect 10275 4981 10284 5015
rect 10232 4972 10284 4981
rect 12900 4972 12952 5024
rect 14556 5015 14608 5024
rect 14556 4981 14565 5015
rect 14565 4981 14599 5015
rect 14599 4981 14608 5015
rect 14556 4972 14608 4981
rect 15936 4972 15988 5024
rect 16764 4972 16816 5024
rect 1918 4870 1970 4922
rect 1982 4870 2034 4922
rect 2046 4870 2098 4922
rect 2110 4870 2162 4922
rect 2174 4870 2226 4922
rect 2238 4870 2290 4922
rect 7918 4870 7970 4922
rect 7982 4870 8034 4922
rect 8046 4870 8098 4922
rect 8110 4870 8162 4922
rect 8174 4870 8226 4922
rect 8238 4870 8290 4922
rect 13918 4870 13970 4922
rect 13982 4870 14034 4922
rect 14046 4870 14098 4922
rect 14110 4870 14162 4922
rect 14174 4870 14226 4922
rect 14238 4870 14290 4922
rect 2320 4811 2372 4820
rect 2320 4777 2329 4811
rect 2329 4777 2363 4811
rect 2363 4777 2372 4811
rect 2320 4768 2372 4777
rect 5448 4768 5500 4820
rect 10048 4768 10100 4820
rect 10692 4768 10744 4820
rect 12256 4768 12308 4820
rect 16580 4768 16632 4820
rect 8392 4700 8444 4752
rect 9128 4700 9180 4752
rect 7564 4632 7616 4684
rect 1584 4607 1636 4616
rect 1584 4573 1593 4607
rect 1593 4573 1627 4607
rect 1627 4573 1636 4607
rect 1584 4564 1636 4573
rect 2412 4607 2464 4616
rect 2412 4573 2421 4607
rect 2421 4573 2455 4607
rect 2455 4573 2464 4607
rect 2412 4564 2464 4573
rect 6368 4607 6420 4616
rect 6368 4573 6377 4607
rect 6377 4573 6411 4607
rect 6411 4573 6420 4607
rect 6368 4564 6420 4573
rect 8576 4564 8628 4616
rect 9312 4675 9364 4684
rect 9312 4641 9321 4675
rect 9321 4641 9355 4675
rect 9355 4641 9364 4675
rect 9312 4632 9364 4641
rect 10508 4700 10560 4752
rect 16672 4743 16724 4752
rect 16672 4709 16681 4743
rect 16681 4709 16715 4743
rect 16715 4709 16724 4743
rect 16672 4700 16724 4709
rect 10876 4632 10928 4684
rect 11152 4675 11204 4684
rect 11152 4641 11161 4675
rect 11161 4641 11195 4675
rect 11195 4641 11204 4675
rect 11152 4632 11204 4641
rect 11612 4632 11664 4684
rect 15568 4632 15620 4684
rect 16028 4632 16080 4684
rect 7196 4496 7248 4548
rect 848 4428 900 4480
rect 6184 4471 6236 4480
rect 6184 4437 6193 4471
rect 6193 4437 6227 4471
rect 6227 4437 6236 4471
rect 6184 4428 6236 4437
rect 7104 4428 7156 4480
rect 7656 4428 7708 4480
rect 9220 4607 9272 4616
rect 9220 4573 9229 4607
rect 9229 4573 9263 4607
rect 9263 4573 9272 4607
rect 9220 4564 9272 4573
rect 9496 4607 9548 4616
rect 9496 4573 9505 4607
rect 9505 4573 9539 4607
rect 9539 4573 9548 4607
rect 9496 4564 9548 4573
rect 10692 4564 10744 4616
rect 11428 4564 11480 4616
rect 16764 4564 16816 4616
rect 13360 4496 13412 4548
rect 13820 4428 13872 4480
rect 2658 4326 2710 4378
rect 2722 4326 2774 4378
rect 2786 4326 2838 4378
rect 2850 4326 2902 4378
rect 2914 4326 2966 4378
rect 2978 4326 3030 4378
rect 8658 4326 8710 4378
rect 8722 4326 8774 4378
rect 8786 4326 8838 4378
rect 8850 4326 8902 4378
rect 8914 4326 8966 4378
rect 8978 4326 9030 4378
rect 14658 4326 14710 4378
rect 14722 4326 14774 4378
rect 14786 4326 14838 4378
rect 14850 4326 14902 4378
rect 14914 4326 14966 4378
rect 14978 4326 15030 4378
rect 4160 4224 4212 4276
rect 8576 4224 8628 4276
rect 10876 4224 10928 4276
rect 11244 4224 11296 4276
rect 11980 4224 12032 4276
rect 12348 4224 12400 4276
rect 12440 4224 12492 4276
rect 13452 4267 13504 4276
rect 13452 4233 13461 4267
rect 13461 4233 13495 4267
rect 13495 4233 13504 4267
rect 13452 4224 13504 4233
rect 14832 4267 14884 4276
rect 14832 4233 14841 4267
rect 14841 4233 14875 4267
rect 14875 4233 14884 4267
rect 14832 4224 14884 4233
rect 11428 4156 11480 4208
rect 3148 4131 3200 4140
rect 3148 4097 3157 4131
rect 3157 4097 3191 4131
rect 3191 4097 3200 4131
rect 3148 4088 3200 4097
rect 3516 4088 3568 4140
rect 1492 4020 1544 4072
rect 6092 4131 6144 4140
rect 6092 4097 6101 4131
rect 6101 4097 6135 4131
rect 6135 4097 6144 4131
rect 6092 4088 6144 4097
rect 6184 4131 6236 4140
rect 6184 4097 6193 4131
rect 6193 4097 6227 4131
rect 6227 4097 6236 4131
rect 6184 4088 6236 4097
rect 6920 4088 6972 4140
rect 4528 3995 4580 4004
rect 4528 3961 4537 3995
rect 4537 3961 4571 3995
rect 4571 3961 4580 3995
rect 4528 3952 4580 3961
rect 5908 3995 5960 4004
rect 5908 3961 5917 3995
rect 5917 3961 5951 3995
rect 5951 3961 5960 3995
rect 5908 3952 5960 3961
rect 6368 4020 6420 4072
rect 7196 4131 7248 4140
rect 7196 4097 7205 4131
rect 7205 4097 7239 4131
rect 7239 4097 7248 4131
rect 7196 4088 7248 4097
rect 7472 4088 7524 4140
rect 8392 4131 8444 4140
rect 8392 4097 8401 4131
rect 8401 4097 8435 4131
rect 8435 4097 8444 4131
rect 8392 4088 8444 4097
rect 9496 4088 9548 4140
rect 6552 3952 6604 4004
rect 6368 3884 6420 3936
rect 8668 4020 8720 4072
rect 7656 3952 7708 4004
rect 10784 3952 10836 4004
rect 12256 4131 12308 4140
rect 12256 4097 12265 4131
rect 12265 4097 12299 4131
rect 12299 4097 12308 4131
rect 12256 4088 12308 4097
rect 12440 4088 12492 4140
rect 12808 4156 12860 4208
rect 13544 4088 13596 4140
rect 14464 4156 14516 4208
rect 15844 4156 15896 4208
rect 13636 4063 13688 4072
rect 13636 4029 13645 4063
rect 13645 4029 13679 4063
rect 13679 4029 13688 4063
rect 13636 4020 13688 4029
rect 12440 3952 12492 4004
rect 14372 4088 14424 4140
rect 15752 4088 15804 4140
rect 11152 3884 11204 3936
rect 11244 3927 11296 3936
rect 11244 3893 11253 3927
rect 11253 3893 11287 3927
rect 11287 3893 11296 3927
rect 11244 3884 11296 3893
rect 12900 3884 12952 3936
rect 13728 3884 13780 3936
rect 15292 4063 15344 4072
rect 15292 4029 15301 4063
rect 15301 4029 15335 4063
rect 15335 4029 15344 4063
rect 15292 4020 15344 4029
rect 15384 4063 15436 4072
rect 15384 4029 15393 4063
rect 15393 4029 15427 4063
rect 15427 4029 15436 4063
rect 15384 4020 15436 4029
rect 15108 3952 15160 4004
rect 14556 3884 14608 3936
rect 15476 3927 15528 3936
rect 15476 3893 15485 3927
rect 15485 3893 15519 3927
rect 15519 3893 15528 3927
rect 15476 3884 15528 3893
rect 1918 3782 1970 3834
rect 1982 3782 2034 3834
rect 2046 3782 2098 3834
rect 2110 3782 2162 3834
rect 2174 3782 2226 3834
rect 2238 3782 2290 3834
rect 7918 3782 7970 3834
rect 7982 3782 8034 3834
rect 8046 3782 8098 3834
rect 8110 3782 8162 3834
rect 8174 3782 8226 3834
rect 8238 3782 8290 3834
rect 13918 3782 13970 3834
rect 13982 3782 14034 3834
rect 14046 3782 14098 3834
rect 14110 3782 14162 3834
rect 14174 3782 14226 3834
rect 14238 3782 14290 3834
rect 4528 3680 4580 3732
rect 8300 3723 8352 3732
rect 8300 3689 8309 3723
rect 8309 3689 8343 3723
rect 8343 3689 8352 3723
rect 8300 3680 8352 3689
rect 6368 3587 6420 3596
rect 6368 3553 6377 3587
rect 6377 3553 6411 3587
rect 6411 3553 6420 3587
rect 6368 3544 6420 3553
rect 6552 3612 6604 3664
rect 8392 3612 8444 3664
rect 10692 3723 10744 3732
rect 10692 3689 10701 3723
rect 10701 3689 10735 3723
rect 10735 3689 10744 3723
rect 10692 3680 10744 3689
rect 12256 3680 12308 3732
rect 13176 3680 13228 3732
rect 13728 3723 13780 3732
rect 13728 3689 13737 3723
rect 13737 3689 13771 3723
rect 13771 3689 13780 3723
rect 13728 3680 13780 3689
rect 14372 3680 14424 3732
rect 14556 3680 14608 3732
rect 12716 3612 12768 3664
rect 12900 3612 12952 3664
rect 13544 3612 13596 3664
rect 14832 3723 14884 3732
rect 14832 3689 14841 3723
rect 14841 3689 14875 3723
rect 14875 3689 14884 3723
rect 14832 3680 14884 3689
rect 15568 3723 15620 3732
rect 15568 3689 15577 3723
rect 15577 3689 15611 3723
rect 15611 3689 15620 3723
rect 15568 3680 15620 3689
rect 3240 3519 3292 3528
rect 3240 3485 3249 3519
rect 3249 3485 3283 3519
rect 3283 3485 3292 3519
rect 3240 3476 3292 3485
rect 6092 3476 6144 3528
rect 4252 3408 4304 3460
rect 848 3340 900 3392
rect 3884 3340 3936 3392
rect 7656 3519 7708 3528
rect 7656 3485 7665 3519
rect 7665 3485 7699 3519
rect 7699 3485 7708 3519
rect 7656 3476 7708 3485
rect 8300 3544 8352 3596
rect 8484 3544 8536 3596
rect 9772 3544 9824 3596
rect 11704 3544 11756 3596
rect 12164 3544 12216 3596
rect 7104 3408 7156 3460
rect 8668 3451 8720 3460
rect 8668 3417 8677 3451
rect 8677 3417 8711 3451
rect 8711 3417 8720 3451
rect 9404 3519 9456 3528
rect 9404 3485 9413 3519
rect 9413 3485 9447 3519
rect 9447 3485 9456 3519
rect 9404 3476 9456 3485
rect 10600 3519 10652 3528
rect 10600 3485 10609 3519
rect 10609 3485 10643 3519
rect 10643 3485 10652 3519
rect 10600 3476 10652 3485
rect 11244 3476 11296 3528
rect 11428 3519 11480 3528
rect 11428 3485 11437 3519
rect 11437 3485 11471 3519
rect 11471 3485 11480 3519
rect 11428 3476 11480 3485
rect 11612 3519 11664 3528
rect 11612 3485 11621 3519
rect 11621 3485 11655 3519
rect 11655 3485 11664 3519
rect 11612 3476 11664 3485
rect 12440 3519 12492 3528
rect 12440 3485 12449 3519
rect 12449 3485 12483 3519
rect 12483 3485 12492 3519
rect 12440 3476 12492 3485
rect 12716 3519 12768 3528
rect 12716 3485 12725 3519
rect 12725 3485 12759 3519
rect 12759 3485 12768 3519
rect 12716 3476 12768 3485
rect 12900 3519 12952 3528
rect 12900 3485 12909 3519
rect 12909 3485 12943 3519
rect 12943 3485 12952 3519
rect 12900 3476 12952 3485
rect 14372 3587 14424 3596
rect 14372 3553 14381 3587
rect 14381 3553 14415 3587
rect 14415 3553 14424 3587
rect 14372 3544 14424 3553
rect 8668 3408 8720 3417
rect 12348 3408 12400 3460
rect 13820 3476 13872 3528
rect 15660 3544 15712 3596
rect 14648 3519 14700 3528
rect 14648 3485 14657 3519
rect 14657 3485 14691 3519
rect 14691 3485 14700 3519
rect 14648 3476 14700 3485
rect 15476 3519 15528 3528
rect 15476 3485 15486 3519
rect 15486 3485 15528 3519
rect 15476 3476 15528 3485
rect 15844 3519 15896 3528
rect 15844 3485 15853 3519
rect 15853 3485 15887 3519
rect 15887 3485 15896 3519
rect 15844 3476 15896 3485
rect 10140 3340 10192 3392
rect 11336 3340 11388 3392
rect 13360 3340 13412 3392
rect 15660 3451 15712 3460
rect 15660 3417 15669 3451
rect 15669 3417 15703 3451
rect 15703 3417 15712 3451
rect 15660 3408 15712 3417
rect 15108 3340 15160 3392
rect 2658 3238 2710 3290
rect 2722 3238 2774 3290
rect 2786 3238 2838 3290
rect 2850 3238 2902 3290
rect 2914 3238 2966 3290
rect 2978 3238 3030 3290
rect 8658 3238 8710 3290
rect 8722 3238 8774 3290
rect 8786 3238 8838 3290
rect 8850 3238 8902 3290
rect 8914 3238 8966 3290
rect 8978 3238 9030 3290
rect 14658 3238 14710 3290
rect 14722 3238 14774 3290
rect 14786 3238 14838 3290
rect 14850 3238 14902 3290
rect 14914 3238 14966 3290
rect 14978 3238 15030 3290
rect 2412 3136 2464 3188
rect 2872 3136 2924 3188
rect 3148 3136 3200 3188
rect 3792 3136 3844 3188
rect 3424 3068 3476 3120
rect 3884 3111 3936 3120
rect 3884 3077 3893 3111
rect 3893 3077 3927 3111
rect 3927 3077 3936 3111
rect 3884 3068 3936 3077
rect 5264 3068 5316 3120
rect 9404 3136 9456 3188
rect 10600 3179 10652 3188
rect 10600 3145 10609 3179
rect 10609 3145 10643 3179
rect 10643 3145 10652 3179
rect 10600 3136 10652 3145
rect 2872 2932 2924 2984
rect 3516 2932 3568 2984
rect 3884 2932 3936 2984
rect 4252 2975 4304 2984
rect 4252 2941 4261 2975
rect 4261 2941 4295 2975
rect 4295 2941 4304 2975
rect 4252 2932 4304 2941
rect 1400 2839 1452 2848
rect 1400 2805 1409 2839
rect 1409 2805 1443 2839
rect 1443 2805 1452 2839
rect 1400 2796 1452 2805
rect 2320 2796 2372 2848
rect 3240 2796 3292 2848
rect 7104 3043 7156 3052
rect 7104 3009 7113 3043
rect 7113 3009 7147 3043
rect 7147 3009 7156 3043
rect 7104 3000 7156 3009
rect 7472 3068 7524 3120
rect 8300 3068 8352 3120
rect 9772 3111 9824 3120
rect 8484 3000 8536 3052
rect 9772 3077 9781 3111
rect 9781 3077 9815 3111
rect 9815 3077 9824 3111
rect 9772 3068 9824 3077
rect 7564 2864 7616 2916
rect 9680 3043 9732 3052
rect 9680 3009 9689 3043
rect 9689 3009 9723 3043
rect 9723 3009 9732 3043
rect 9680 3000 9732 3009
rect 10140 3043 10192 3052
rect 10140 3009 10149 3043
rect 10149 3009 10183 3043
rect 10183 3009 10192 3043
rect 10876 3068 10928 3120
rect 11704 3179 11756 3188
rect 11704 3145 11713 3179
rect 11713 3145 11747 3179
rect 11747 3145 11756 3179
rect 11704 3136 11756 3145
rect 12348 3136 12400 3188
rect 14556 3136 14608 3188
rect 15108 3179 15160 3188
rect 15108 3145 15117 3179
rect 15117 3145 15151 3179
rect 15151 3145 15160 3179
rect 15108 3136 15160 3145
rect 10140 3000 10192 3009
rect 11152 3068 11204 3120
rect 12716 3068 12768 3120
rect 13544 3068 13596 3120
rect 10876 2932 10928 2984
rect 11980 3043 12032 3052
rect 11980 3009 11989 3043
rect 11989 3009 12023 3043
rect 12023 3009 12032 3043
rect 11980 3000 12032 3009
rect 11060 2864 11112 2916
rect 10784 2839 10836 2848
rect 10784 2805 10793 2839
rect 10793 2805 10827 2839
rect 10827 2805 10836 2839
rect 10784 2796 10836 2805
rect 10876 2796 10928 2848
rect 12440 3000 12492 3052
rect 13728 3000 13780 3052
rect 15752 3068 15804 3120
rect 15568 3000 15620 3052
rect 11980 2864 12032 2916
rect 12900 2932 12952 2984
rect 14372 2907 14424 2916
rect 12348 2796 12400 2848
rect 14372 2873 14381 2907
rect 14381 2873 14415 2907
rect 14415 2873 14424 2907
rect 14372 2864 14424 2873
rect 15660 2864 15712 2916
rect 12716 2796 12768 2848
rect 13636 2796 13688 2848
rect 1918 2694 1970 2746
rect 1982 2694 2034 2746
rect 2046 2694 2098 2746
rect 2110 2694 2162 2746
rect 2174 2694 2226 2746
rect 2238 2694 2290 2746
rect 7918 2694 7970 2746
rect 7982 2694 8034 2746
rect 8046 2694 8098 2746
rect 8110 2694 8162 2746
rect 8174 2694 8226 2746
rect 8238 2694 8290 2746
rect 13918 2694 13970 2746
rect 13982 2694 14034 2746
rect 14046 2694 14098 2746
rect 14110 2694 14162 2746
rect 14174 2694 14226 2746
rect 14238 2694 14290 2746
rect 1584 2592 1636 2644
rect 3424 2592 3476 2644
rect 5264 2592 5316 2644
rect 9680 2592 9732 2644
rect 13176 2635 13228 2644
rect 13176 2601 13185 2635
rect 13185 2601 13219 2635
rect 13219 2601 13228 2635
rect 13176 2592 13228 2601
rect 12900 2524 12952 2576
rect 3792 2456 3844 2508
rect 3976 2431 4028 2440
rect 3976 2397 3985 2431
rect 3985 2397 4019 2431
rect 4019 2397 4028 2431
rect 3976 2388 4028 2397
rect 12992 2456 13044 2508
rect 9404 2388 9456 2440
rect 11428 2388 11480 2440
rect 12348 2388 12400 2440
rect 12716 2388 12768 2440
rect 2320 2320 2372 2372
rect 7564 2320 7616 2372
rect 2658 2150 2710 2202
rect 2722 2150 2774 2202
rect 2786 2150 2838 2202
rect 2850 2150 2902 2202
rect 2914 2150 2966 2202
rect 2978 2150 3030 2202
rect 8658 2150 8710 2202
rect 8722 2150 8774 2202
rect 8786 2150 8838 2202
rect 8850 2150 8902 2202
rect 8914 2150 8966 2202
rect 8978 2150 9030 2202
rect 14658 2150 14710 2202
rect 14722 2150 14774 2202
rect 14786 2150 14838 2202
rect 14850 2150 14902 2202
rect 14914 2150 14966 2202
rect 14978 2150 15030 2202
<< metal2 >>
rect 1122 20301 1178 21101
rect 2226 20301 2282 21101
rect 3330 20301 3386 21101
rect 4434 20301 4490 21101
rect 5538 20301 5594 21101
rect 6642 20301 6698 21101
rect 7746 20301 7802 21101
rect 8850 20301 8906 21101
rect 8956 20318 9168 20346
rect 1136 18290 1164 20301
rect 1214 18592 1270 18601
rect 1214 18527 1270 18536
rect 1228 18426 1256 18527
rect 1216 18420 1268 18426
rect 1216 18362 1268 18368
rect 2240 18290 2268 20301
rect 2656 18524 3032 18533
rect 2712 18522 2736 18524
rect 2792 18522 2816 18524
rect 2872 18522 2896 18524
rect 2952 18522 2976 18524
rect 2712 18470 2722 18522
rect 2966 18470 2976 18522
rect 2712 18468 2736 18470
rect 2792 18468 2816 18470
rect 2872 18468 2896 18470
rect 2952 18468 2976 18470
rect 2656 18459 3032 18468
rect 3344 18290 3372 20301
rect 4448 18290 4476 20301
rect 5552 18290 5580 20301
rect 5724 18420 5776 18426
rect 5724 18362 5776 18368
rect 1124 18284 1176 18290
rect 1124 18226 1176 18232
rect 2228 18284 2280 18290
rect 2228 18226 2280 18232
rect 3332 18284 3384 18290
rect 3332 18226 3384 18232
rect 4436 18284 4488 18290
rect 4436 18226 4488 18232
rect 5540 18284 5592 18290
rect 5540 18226 5592 18232
rect 3516 18216 3568 18222
rect 3516 18158 3568 18164
rect 1584 18080 1636 18086
rect 1584 18022 1636 18028
rect 1596 17610 1624 18022
rect 1916 17980 2292 17989
rect 1972 17978 1996 17980
rect 2052 17978 2076 17980
rect 2132 17978 2156 17980
rect 2212 17978 2236 17980
rect 1972 17926 1982 17978
rect 2226 17926 2236 17978
rect 1972 17924 1996 17926
rect 2052 17924 2076 17926
rect 2132 17924 2156 17926
rect 2212 17924 2236 17926
rect 1916 17915 2292 17924
rect 1584 17604 1636 17610
rect 1584 17546 1636 17552
rect 2228 17604 2280 17610
rect 2228 17546 2280 17552
rect 3240 17604 3292 17610
rect 3240 17546 3292 17552
rect 1306 17504 1362 17513
rect 1306 17439 1362 17448
rect 1320 17338 1348 17439
rect 2240 17338 2268 17546
rect 2504 17536 2556 17542
rect 2504 17478 2556 17484
rect 1308 17332 1360 17338
rect 1308 17274 1360 17280
rect 2228 17332 2280 17338
rect 2228 17274 2280 17280
rect 2516 17202 2544 17478
rect 2656 17436 3032 17445
rect 2712 17434 2736 17436
rect 2792 17434 2816 17436
rect 2872 17434 2896 17436
rect 2952 17434 2976 17436
rect 2712 17382 2722 17434
rect 2966 17382 2976 17434
rect 2712 17380 2736 17382
rect 2792 17380 2816 17382
rect 2872 17380 2896 17382
rect 2952 17380 2976 17382
rect 2656 17371 3032 17380
rect 2504 17196 2556 17202
rect 2504 17138 2556 17144
rect 1916 16892 2292 16901
rect 1972 16890 1996 16892
rect 2052 16890 2076 16892
rect 2132 16890 2156 16892
rect 2212 16890 2236 16892
rect 1972 16838 1982 16890
rect 2226 16838 2236 16890
rect 1972 16836 1996 16838
rect 2052 16836 2076 16838
rect 2132 16836 2156 16838
rect 2212 16836 2236 16838
rect 1916 16827 2292 16836
rect 1400 16584 1452 16590
rect 846 16552 902 16561
rect 1400 16526 1452 16532
rect 846 16487 902 16496
rect 860 16454 888 16487
rect 848 16448 900 16454
rect 848 16390 900 16396
rect 848 15904 900 15910
rect 848 15846 900 15852
rect 860 15473 888 15846
rect 1412 15706 1440 16526
rect 2516 16114 2544 17138
rect 3056 17128 3108 17134
rect 3056 17070 3108 17076
rect 2656 16348 3032 16357
rect 2712 16346 2736 16348
rect 2792 16346 2816 16348
rect 2872 16346 2896 16348
rect 2952 16346 2976 16348
rect 2712 16294 2722 16346
rect 2966 16294 2976 16346
rect 2712 16292 2736 16294
rect 2792 16292 2816 16294
rect 2872 16292 2896 16294
rect 2952 16292 2976 16294
rect 2656 16283 3032 16292
rect 3068 16250 3096 17070
rect 3056 16244 3108 16250
rect 3056 16186 3108 16192
rect 1584 16108 1636 16114
rect 1584 16050 1636 16056
rect 2504 16108 2556 16114
rect 2504 16050 2556 16056
rect 1400 15700 1452 15706
rect 1400 15642 1452 15648
rect 846 15464 902 15473
rect 846 15399 902 15408
rect 1596 15162 1624 16050
rect 2320 15904 2372 15910
rect 2320 15846 2372 15852
rect 1916 15804 2292 15813
rect 1972 15802 1996 15804
rect 2052 15802 2076 15804
rect 2132 15802 2156 15804
rect 2212 15802 2236 15804
rect 1972 15750 1982 15802
rect 2226 15750 2236 15802
rect 1972 15748 1996 15750
rect 2052 15748 2076 15750
rect 2132 15748 2156 15750
rect 2212 15748 2236 15750
rect 1916 15739 2292 15748
rect 2332 15434 2360 15846
rect 2320 15428 2372 15434
rect 2320 15370 2372 15376
rect 1584 15156 1636 15162
rect 1584 15098 1636 15104
rect 2412 15088 2464 15094
rect 2412 15030 2464 15036
rect 1916 14716 2292 14725
rect 1972 14714 1996 14716
rect 2052 14714 2076 14716
rect 2132 14714 2156 14716
rect 2212 14714 2236 14716
rect 1972 14662 1982 14714
rect 2226 14662 2236 14714
rect 1972 14660 1996 14662
rect 2052 14660 2076 14662
rect 2132 14660 2156 14662
rect 2212 14660 2236 14662
rect 1916 14651 2292 14660
rect 2424 14618 2452 15030
rect 2412 14612 2464 14618
rect 2412 14554 2464 14560
rect 2516 14414 2544 16050
rect 3148 16040 3200 16046
rect 3148 15982 3200 15988
rect 3160 15502 3188 15982
rect 3148 15496 3200 15502
rect 3148 15438 3200 15444
rect 2656 15260 3032 15269
rect 2712 15258 2736 15260
rect 2792 15258 2816 15260
rect 2872 15258 2896 15260
rect 2952 15258 2976 15260
rect 2712 15206 2722 15258
rect 2966 15206 2976 15258
rect 2712 15204 2736 15206
rect 2792 15204 2816 15206
rect 2872 15204 2896 15206
rect 2952 15204 2976 15206
rect 2656 15195 3032 15204
rect 3160 14958 3188 15438
rect 2872 14952 2924 14958
rect 2872 14894 2924 14900
rect 3148 14952 3200 14958
rect 3252 14929 3280 17546
rect 3528 17338 3556 18158
rect 4896 18080 4948 18086
rect 4896 18022 4948 18028
rect 4068 17740 4120 17746
rect 4068 17682 4120 17688
rect 4080 17626 4108 17682
rect 3988 17598 4108 17626
rect 4908 17610 4936 18022
rect 4896 17604 4948 17610
rect 3884 17536 3936 17542
rect 3884 17478 3936 17484
rect 3516 17332 3568 17338
rect 3516 17274 3568 17280
rect 3332 16652 3384 16658
rect 3332 16594 3384 16600
rect 3344 15706 3372 16594
rect 3896 16182 3924 17478
rect 3988 16998 4016 17598
rect 4896 17546 4948 17552
rect 4436 17536 4488 17542
rect 4436 17478 4488 17484
rect 4448 17270 4476 17478
rect 4436 17264 4488 17270
rect 4436 17206 4488 17212
rect 4252 17128 4304 17134
rect 4252 17070 4304 17076
rect 3976 16992 4028 16998
rect 3976 16934 4028 16940
rect 3884 16176 3936 16182
rect 3884 16118 3936 16124
rect 3988 16046 4016 16934
rect 4068 16584 4120 16590
rect 4068 16526 4120 16532
rect 4080 16250 4108 16526
rect 4160 16448 4212 16454
rect 4264 16436 4292 17070
rect 4344 16788 4396 16794
rect 4344 16730 4396 16736
rect 4212 16408 4292 16436
rect 4160 16390 4212 16396
rect 4068 16244 4120 16250
rect 4068 16186 4120 16192
rect 4356 16182 4384 16730
rect 4344 16176 4396 16182
rect 4344 16118 4396 16124
rect 3976 16040 4028 16046
rect 3976 15982 4028 15988
rect 3332 15700 3384 15706
rect 3332 15642 3384 15648
rect 4252 15564 4304 15570
rect 4252 15506 4304 15512
rect 4264 15162 4292 15506
rect 4252 15156 4304 15162
rect 4252 15098 4304 15104
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 3148 14894 3200 14900
rect 3238 14920 3294 14929
rect 2884 14618 2912 14894
rect 2872 14612 2924 14618
rect 2872 14554 2924 14560
rect 1400 14408 1452 14414
rect 846 14376 902 14385
rect 1400 14350 1452 14356
rect 2504 14408 2556 14414
rect 2504 14350 2556 14356
rect 846 14311 902 14320
rect 860 14278 888 14311
rect 848 14272 900 14278
rect 848 14214 900 14220
rect 1412 14074 1440 14350
rect 1400 14068 1452 14074
rect 1400 14010 1452 14016
rect 2320 14000 2372 14006
rect 2320 13942 2372 13948
rect 1916 13628 2292 13637
rect 1972 13626 1996 13628
rect 2052 13626 2076 13628
rect 2132 13626 2156 13628
rect 2212 13626 2236 13628
rect 1972 13574 1982 13626
rect 2226 13574 2236 13626
rect 1972 13572 1996 13574
rect 2052 13572 2076 13574
rect 2132 13572 2156 13574
rect 2212 13572 2236 13574
rect 1916 13563 2292 13572
rect 2332 13530 2360 13942
rect 2320 13524 2372 13530
rect 2320 13466 2372 13472
rect 2516 13326 2544 14350
rect 2656 14172 3032 14181
rect 2712 14170 2736 14172
rect 2792 14170 2816 14172
rect 2872 14170 2896 14172
rect 2952 14170 2976 14172
rect 2712 14118 2722 14170
rect 2966 14118 2976 14170
rect 2712 14116 2736 14118
rect 2792 14116 2816 14118
rect 2872 14116 2896 14118
rect 2952 14116 2976 14118
rect 2656 14107 3032 14116
rect 3160 13870 3188 14894
rect 3238 14855 3294 14864
rect 2872 13864 2924 13870
rect 2872 13806 2924 13812
rect 3148 13864 3200 13870
rect 3148 13806 3200 13812
rect 2884 13530 2912 13806
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 1400 13320 1452 13326
rect 846 13288 902 13297
rect 1400 13262 1452 13268
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 846 13223 902 13232
rect 860 13190 888 13223
rect 848 13184 900 13190
rect 848 13126 900 13132
rect 1412 12986 1440 13262
rect 1400 12980 1452 12986
rect 1400 12922 1452 12928
rect 2320 12912 2372 12918
rect 2320 12854 2372 12860
rect 1916 12540 2292 12549
rect 1972 12538 1996 12540
rect 2052 12538 2076 12540
rect 2132 12538 2156 12540
rect 2212 12538 2236 12540
rect 1972 12486 1982 12538
rect 2226 12486 2236 12538
rect 1972 12484 1996 12486
rect 2052 12484 2076 12486
rect 2132 12484 2156 12486
rect 2212 12484 2236 12486
rect 1916 12475 2292 12484
rect 2332 12442 2360 12854
rect 2320 12436 2372 12442
rect 2320 12378 2372 12384
rect 2516 12238 2544 13262
rect 2656 13084 3032 13093
rect 2712 13082 2736 13084
rect 2792 13082 2816 13084
rect 2872 13082 2896 13084
rect 2952 13082 2976 13084
rect 2712 13030 2722 13082
rect 2966 13030 2976 13082
rect 2712 13028 2736 13030
rect 2792 13028 2816 13030
rect 2872 13028 2896 13030
rect 2952 13028 2976 13030
rect 2656 13019 3032 13028
rect 3160 12646 3188 13806
rect 3148 12640 3200 12646
rect 3148 12582 3200 12588
rect 1400 12232 1452 12238
rect 846 12200 902 12209
rect 1400 12174 1452 12180
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 846 12135 902 12144
rect 860 12102 888 12135
rect 848 12096 900 12102
rect 848 12038 900 12044
rect 1412 11354 1440 12174
rect 1916 11452 2292 11461
rect 1972 11450 1996 11452
rect 2052 11450 2076 11452
rect 2132 11450 2156 11452
rect 2212 11450 2236 11452
rect 1972 11398 1982 11450
rect 2226 11398 2236 11450
rect 1972 11396 1996 11398
rect 2052 11396 2076 11398
rect 2132 11396 2156 11398
rect 2212 11396 2236 11398
rect 1916 11387 2292 11396
rect 1400 11348 1452 11354
rect 1400 11290 1452 11296
rect 2516 11014 2544 12174
rect 2656 11996 3032 12005
rect 2712 11994 2736 11996
rect 2792 11994 2816 11996
rect 2872 11994 2896 11996
rect 2952 11994 2976 11996
rect 2712 11942 2722 11994
rect 2966 11942 2976 11994
rect 2712 11940 2736 11942
rect 2792 11940 2816 11942
rect 2872 11940 2896 11942
rect 2952 11940 2976 11942
rect 2656 11931 3032 11940
rect 3160 11218 3188 12582
rect 3148 11212 3200 11218
rect 3148 11154 3200 11160
rect 2504 11008 2556 11014
rect 1306 10976 1362 10985
rect 2504 10950 2556 10956
rect 1306 10911 1362 10920
rect 1320 10810 1348 10911
rect 1308 10804 1360 10810
rect 1308 10746 1360 10752
rect 1400 10668 1452 10674
rect 1400 10610 1452 10616
rect 1412 10266 1440 10610
rect 1916 10364 2292 10373
rect 1972 10362 1996 10364
rect 2052 10362 2076 10364
rect 2132 10362 2156 10364
rect 2212 10362 2236 10364
rect 1972 10310 1982 10362
rect 2226 10310 2236 10362
rect 1972 10308 1996 10310
rect 2052 10308 2076 10310
rect 2132 10308 2156 10310
rect 2212 10308 2236 10310
rect 1916 10299 2292 10308
rect 1400 10260 1452 10266
rect 1400 10202 1452 10208
rect 2412 9988 2464 9994
rect 2412 9930 2464 9936
rect 1306 9888 1362 9897
rect 1306 9823 1362 9832
rect 1320 9450 1348 9823
rect 2424 9654 2452 9930
rect 2516 9926 2544 10950
rect 2656 10908 3032 10917
rect 2712 10906 2736 10908
rect 2792 10906 2816 10908
rect 2872 10906 2896 10908
rect 2952 10906 2976 10908
rect 2712 10854 2722 10906
rect 2966 10854 2976 10906
rect 2712 10852 2736 10854
rect 2792 10852 2816 10854
rect 2872 10852 2896 10854
rect 2952 10852 2976 10854
rect 2656 10843 3032 10852
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 2504 9920 2556 9926
rect 2504 9862 2556 9868
rect 2412 9648 2464 9654
rect 2412 9590 2464 9596
rect 2516 9586 2544 9862
rect 2656 9820 3032 9829
rect 2712 9818 2736 9820
rect 2792 9818 2816 9820
rect 2872 9818 2896 9820
rect 2952 9818 2976 9820
rect 2712 9766 2722 9818
rect 2966 9766 2976 9818
rect 2712 9764 2736 9766
rect 2792 9764 2816 9766
rect 2872 9764 2896 9766
rect 2952 9764 2976 9766
rect 2656 9755 3032 9764
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 2504 9580 2556 9586
rect 2504 9522 2556 9528
rect 1308 9444 1360 9450
rect 1308 9386 1360 9392
rect 1412 9178 1440 9522
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 1916 9276 2292 9285
rect 1972 9274 1996 9276
rect 2052 9274 2076 9276
rect 2132 9274 2156 9276
rect 2212 9274 2236 9276
rect 1972 9222 1982 9274
rect 2226 9222 2236 9274
rect 1972 9220 1996 9222
rect 2052 9220 2076 9222
rect 2132 9220 2156 9222
rect 2212 9220 2236 9222
rect 1916 9211 2292 9220
rect 1400 9172 1452 9178
rect 1400 9114 1452 9120
rect 2228 8900 2280 8906
rect 2228 8842 2280 8848
rect 1306 8800 1362 8809
rect 1306 8735 1362 8744
rect 1320 8634 1348 8735
rect 2240 8634 2268 8842
rect 1308 8628 1360 8634
rect 1308 8570 1360 8576
rect 2228 8628 2280 8634
rect 2228 8570 2280 8576
rect 2424 8498 2452 9454
rect 3160 9450 3188 9998
rect 3148 9444 3200 9450
rect 3148 9386 3200 9392
rect 3160 9042 3188 9386
rect 3148 9036 3200 9042
rect 3148 8978 3200 8984
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 2656 8732 3032 8741
rect 2712 8730 2736 8732
rect 2792 8730 2816 8732
rect 2872 8730 2896 8732
rect 2952 8730 2976 8732
rect 2712 8678 2722 8730
rect 2966 8678 2976 8730
rect 2712 8676 2736 8678
rect 2792 8676 2816 8678
rect 2872 8676 2896 8678
rect 2952 8676 2976 8678
rect 2656 8667 3032 8676
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 2412 8492 2464 8498
rect 2412 8434 2464 8440
rect 1596 8090 1624 8434
rect 1916 8188 2292 8197
rect 1972 8186 1996 8188
rect 2052 8186 2076 8188
rect 2132 8186 2156 8188
rect 2212 8186 2236 8188
rect 1972 8134 1982 8186
rect 2226 8134 2236 8186
rect 1972 8132 1996 8134
rect 2052 8132 2076 8134
rect 2132 8132 2156 8134
rect 2212 8132 2236 8134
rect 1916 8123 2292 8132
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 2320 7812 2372 7818
rect 2320 7754 2372 7760
rect 1306 7712 1362 7721
rect 1306 7647 1362 7656
rect 1320 7546 1348 7647
rect 2332 7546 2360 7754
rect 1308 7540 1360 7546
rect 1308 7482 1360 7488
rect 2320 7540 2372 7546
rect 2320 7482 2372 7488
rect 2424 7410 2452 8434
rect 3068 8430 3096 8774
rect 3056 8424 3108 8430
rect 3056 8366 3108 8372
rect 3160 7954 3188 8978
rect 3148 7948 3200 7954
rect 3148 7890 3200 7896
rect 2656 7644 3032 7653
rect 2712 7642 2736 7644
rect 2792 7642 2816 7644
rect 2872 7642 2896 7644
rect 2952 7642 2976 7644
rect 2712 7590 2722 7642
rect 2966 7590 2976 7642
rect 2712 7588 2736 7590
rect 2792 7588 2816 7590
rect 2872 7588 2896 7590
rect 2952 7588 2976 7590
rect 2656 7579 3032 7588
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 2412 7404 2464 7410
rect 2412 7346 2464 7352
rect 1596 7002 1624 7346
rect 1916 7100 2292 7109
rect 1972 7098 1996 7100
rect 2052 7098 2076 7100
rect 2132 7098 2156 7100
rect 2212 7098 2236 7100
rect 1972 7046 1982 7098
rect 2226 7046 2236 7098
rect 1972 7044 1996 7046
rect 2052 7044 2076 7046
rect 2132 7044 2156 7046
rect 2212 7044 2236 7046
rect 1916 7035 2292 7044
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 2320 6724 2372 6730
rect 2320 6666 2372 6672
rect 1306 6624 1362 6633
rect 1306 6559 1362 6568
rect 1320 6458 1348 6559
rect 2332 6458 2360 6666
rect 1308 6452 1360 6458
rect 1308 6394 1360 6400
rect 2320 6452 2372 6458
rect 2320 6394 2372 6400
rect 2424 6322 2452 7346
rect 3160 6866 3188 7890
rect 3148 6860 3200 6866
rect 3148 6802 3200 6808
rect 2656 6556 3032 6565
rect 2712 6554 2736 6556
rect 2792 6554 2816 6556
rect 2872 6554 2896 6556
rect 2952 6554 2976 6556
rect 2712 6502 2722 6554
rect 2966 6502 2976 6554
rect 2712 6500 2736 6502
rect 2792 6500 2816 6502
rect 2872 6500 2896 6502
rect 2952 6500 2976 6502
rect 2656 6491 3032 6500
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 1492 5704 1544 5710
rect 1492 5646 1544 5652
rect 1400 5568 1452 5574
rect 1398 5536 1400 5545
rect 1452 5536 1454 5545
rect 1398 5471 1454 5480
rect 846 4584 902 4593
rect 846 4519 902 4528
rect 860 4486 888 4519
rect 848 4480 900 4486
rect 848 4422 900 4428
rect 1504 4078 1532 5646
rect 1596 5370 1624 6258
rect 1916 6012 2292 6021
rect 1972 6010 1996 6012
rect 2052 6010 2076 6012
rect 2132 6010 2156 6012
rect 2212 6010 2236 6012
rect 1972 5958 1982 6010
rect 2226 5958 2236 6010
rect 1972 5956 1996 5958
rect 2052 5956 2076 5958
rect 2132 5956 2156 5958
rect 2212 5956 2236 5958
rect 1916 5947 2292 5956
rect 1584 5364 1636 5370
rect 1584 5306 1636 5312
rect 2320 5296 2372 5302
rect 2320 5238 2372 5244
rect 1916 4924 2292 4933
rect 1972 4922 1996 4924
rect 2052 4922 2076 4924
rect 2132 4922 2156 4924
rect 2212 4922 2236 4924
rect 1972 4870 1982 4922
rect 2226 4870 2236 4922
rect 1972 4868 1996 4870
rect 2052 4868 2076 4870
rect 2132 4868 2156 4870
rect 2212 4868 2236 4870
rect 1916 4859 2292 4868
rect 2332 4826 2360 5238
rect 2320 4820 2372 4826
rect 2320 4762 2372 4768
rect 2424 4622 2452 6258
rect 2656 5468 3032 5477
rect 2712 5466 2736 5468
rect 2792 5466 2816 5468
rect 2872 5466 2896 5468
rect 2952 5466 2976 5468
rect 2712 5414 2722 5466
rect 2966 5414 2976 5466
rect 2712 5412 2736 5414
rect 2792 5412 2816 5414
rect 2872 5412 2896 5414
rect 2952 5412 2976 5414
rect 2656 5403 3032 5412
rect 3160 5234 3188 6802
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 1492 4072 1544 4078
rect 1492 4014 1544 4020
rect 846 3496 902 3505
rect 846 3431 902 3440
rect 860 3398 888 3431
rect 848 3392 900 3398
rect 848 3334 900 3340
rect 1400 2848 1452 2854
rect 1400 2790 1452 2796
rect 1412 2281 1440 2790
rect 1596 2650 1624 4558
rect 1916 3836 2292 3845
rect 1972 3834 1996 3836
rect 2052 3834 2076 3836
rect 2132 3834 2156 3836
rect 2212 3834 2236 3836
rect 1972 3782 1982 3834
rect 2226 3782 2236 3834
rect 1972 3780 1996 3782
rect 2052 3780 2076 3782
rect 2132 3780 2156 3782
rect 2212 3780 2236 3782
rect 1916 3771 2292 3780
rect 2424 3194 2452 4558
rect 2656 4380 3032 4389
rect 2712 4378 2736 4380
rect 2792 4378 2816 4380
rect 2872 4378 2896 4380
rect 2952 4378 2976 4380
rect 2712 4326 2722 4378
rect 2966 4326 2976 4378
rect 2712 4324 2736 4326
rect 2792 4324 2816 4326
rect 2872 4324 2896 4326
rect 2952 4324 2976 4326
rect 2656 4315 3032 4324
rect 3160 4146 3188 5170
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 2656 3292 3032 3301
rect 2712 3290 2736 3292
rect 2792 3290 2816 3292
rect 2872 3290 2896 3292
rect 2952 3290 2976 3292
rect 2712 3238 2722 3290
rect 2966 3238 2976 3290
rect 2712 3236 2736 3238
rect 2792 3236 2816 3238
rect 2872 3236 2896 3238
rect 2952 3236 2976 3238
rect 2656 3227 3032 3236
rect 3160 3194 3188 4082
rect 3252 3534 3280 14855
rect 4080 14600 4108 14962
rect 4436 14952 4488 14958
rect 4436 14894 4488 14900
rect 4620 14952 4672 14958
rect 4620 14894 4672 14900
rect 5356 14952 5408 14958
rect 5356 14894 5408 14900
rect 4344 14612 4396 14618
rect 4080 14572 4344 14600
rect 4080 14346 4108 14572
rect 4344 14554 4396 14560
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 4068 14340 4120 14346
rect 4068 14282 4120 14288
rect 3516 13320 3568 13326
rect 3516 13262 3568 13268
rect 3528 12986 3556 13262
rect 3516 12980 3568 12986
rect 3516 12922 3568 12928
rect 3424 12844 3476 12850
rect 3424 12786 3476 12792
rect 3436 12442 3464 12786
rect 3608 12708 3660 12714
rect 3608 12650 3660 12656
rect 3424 12436 3476 12442
rect 3424 12378 3476 12384
rect 3436 11762 3464 12378
rect 3620 11898 3648 12650
rect 4080 12442 4108 14282
rect 4172 14278 4200 14350
rect 4448 14346 4476 14894
rect 4632 14346 4660 14894
rect 5368 14618 5396 14894
rect 5356 14612 5408 14618
rect 5356 14554 5408 14560
rect 5368 14414 5396 14554
rect 4988 14408 5040 14414
rect 4988 14350 5040 14356
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 4436 14340 4488 14346
rect 4436 14282 4488 14288
rect 4620 14340 4672 14346
rect 4620 14282 4672 14288
rect 4160 14272 4212 14278
rect 4160 14214 4212 14220
rect 5000 13190 5028 14350
rect 5264 13524 5316 13530
rect 5264 13466 5316 13472
rect 5276 13326 5304 13466
rect 5356 13388 5408 13394
rect 5356 13330 5408 13336
rect 5264 13320 5316 13326
rect 5264 13262 5316 13268
rect 4988 13184 5040 13190
rect 4988 13126 5040 13132
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 5172 12844 5224 12850
rect 5276 12832 5304 13262
rect 5368 12986 5396 13330
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 5356 12844 5408 12850
rect 5276 12804 5356 12832
rect 5172 12786 5224 12792
rect 5540 12844 5592 12850
rect 5356 12786 5408 12792
rect 5460 12804 5540 12832
rect 4252 12708 4304 12714
rect 4252 12650 4304 12656
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 4264 12374 4292 12650
rect 4724 12442 4752 12786
rect 4988 12776 5040 12782
rect 4988 12718 5040 12724
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 4252 12368 4304 12374
rect 4252 12310 4304 12316
rect 4160 12232 4212 12238
rect 4160 12174 4212 12180
rect 3700 12164 3752 12170
rect 3700 12106 3752 12112
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 3712 11626 3740 12106
rect 4172 11762 4200 12174
rect 4160 11756 4212 11762
rect 4160 11698 4212 11704
rect 4264 11694 4292 12310
rect 5000 12306 5028 12718
rect 5184 12374 5212 12786
rect 5172 12368 5224 12374
rect 5172 12310 5224 12316
rect 4988 12300 5040 12306
rect 4988 12242 5040 12248
rect 4528 12232 4580 12238
rect 4528 12174 4580 12180
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 4356 11898 4384 12038
rect 4344 11892 4396 11898
rect 4344 11834 4396 11840
rect 4540 11762 4568 12174
rect 5460 11898 5488 12804
rect 5540 12786 5592 12792
rect 5644 12714 5672 13262
rect 5632 12708 5684 12714
rect 5632 12650 5684 12656
rect 5644 12442 5672 12650
rect 5632 12436 5684 12442
rect 5632 12378 5684 12384
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 4528 11756 4580 11762
rect 4528 11698 4580 11704
rect 4804 11756 4856 11762
rect 4804 11698 4856 11704
rect 4252 11688 4304 11694
rect 4252 11630 4304 11636
rect 3700 11620 3752 11626
rect 3700 11562 3752 11568
rect 3712 11218 3740 11562
rect 4816 11354 4844 11698
rect 5460 11354 5488 11834
rect 4804 11348 4856 11354
rect 4804 11290 4856 11296
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 3700 11212 3752 11218
rect 3700 11154 3752 11160
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 3436 9382 3464 9522
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3436 8430 3464 9318
rect 3528 9178 3556 9522
rect 3712 9518 3740 11154
rect 5736 10606 5764 18362
rect 6656 18358 6684 20301
rect 7760 19122 7788 20301
rect 8864 20210 8892 20301
rect 8956 20210 8984 20318
rect 8864 20182 8984 20210
rect 7760 19094 7972 19122
rect 7012 18420 7064 18426
rect 7012 18362 7064 18368
rect 6644 18352 6696 18358
rect 6644 18294 6696 18300
rect 6368 18216 6420 18222
rect 6368 18158 6420 18164
rect 6380 17746 6408 18158
rect 7024 17746 7052 18362
rect 7104 18352 7156 18358
rect 7104 18294 7156 18300
rect 6368 17740 6420 17746
rect 6368 17682 6420 17688
rect 7012 17740 7064 17746
rect 7012 17682 7064 17688
rect 6460 17604 6512 17610
rect 6460 17546 6512 17552
rect 6644 17604 6696 17610
rect 6644 17546 6696 17552
rect 6472 17338 6500 17546
rect 6552 17536 6604 17542
rect 6552 17478 6604 17484
rect 6460 17332 6512 17338
rect 6460 17274 6512 17280
rect 6564 17202 6592 17478
rect 6552 17196 6604 17202
rect 6552 17138 6604 17144
rect 5816 16652 5868 16658
rect 5816 16594 5868 16600
rect 5828 16250 5856 16594
rect 6552 16448 6604 16454
rect 6552 16390 6604 16396
rect 5816 16244 5868 16250
rect 5816 16186 5868 16192
rect 6564 16114 6592 16390
rect 6552 16108 6604 16114
rect 6552 16050 6604 16056
rect 6092 14816 6144 14822
rect 6092 14758 6144 14764
rect 6104 14550 6132 14758
rect 6092 14544 6144 14550
rect 6092 14486 6144 14492
rect 6104 14414 6132 14486
rect 6092 14408 6144 14414
rect 6092 14350 6144 14356
rect 6368 13728 6420 13734
rect 6368 13670 6420 13676
rect 6380 13326 6408 13670
rect 6368 13320 6420 13326
rect 6368 13262 6420 13268
rect 6368 13184 6420 13190
rect 6368 13126 6420 13132
rect 6380 12782 6408 13126
rect 6368 12776 6420 12782
rect 6368 12718 6420 12724
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 6196 11898 6224 12174
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 6380 10674 6408 12718
rect 6656 12102 6684 17546
rect 7116 17338 7144 18294
rect 7944 18290 7972 19094
rect 8656 18524 9032 18533
rect 8712 18522 8736 18524
rect 8792 18522 8816 18524
rect 8872 18522 8896 18524
rect 8952 18522 8976 18524
rect 8712 18470 8722 18522
rect 8966 18470 8976 18522
rect 8712 18468 8736 18470
rect 8792 18468 8816 18470
rect 8872 18468 8896 18470
rect 8952 18468 8976 18470
rect 8656 18459 9032 18468
rect 9140 18290 9168 20318
rect 9954 20301 10010 21101
rect 11058 20301 11114 21101
rect 12162 20301 12218 21101
rect 13266 20301 13322 21101
rect 14370 20301 14426 21101
rect 15474 20301 15530 21101
rect 16578 20301 16634 21101
rect 17682 20301 17738 21101
rect 9968 18290 9996 20301
rect 11072 19258 11100 20301
rect 11072 19230 11192 19258
rect 11164 18290 11192 19230
rect 12176 18290 12204 20301
rect 13280 18290 13308 20301
rect 14384 18290 14412 20301
rect 14656 18524 15032 18533
rect 14712 18522 14736 18524
rect 14792 18522 14816 18524
rect 14872 18522 14896 18524
rect 14952 18522 14976 18524
rect 14712 18470 14722 18522
rect 14966 18470 14976 18522
rect 14712 18468 14736 18470
rect 14792 18468 14816 18470
rect 14872 18468 14896 18470
rect 14952 18468 14976 18470
rect 14656 18459 15032 18468
rect 15488 18290 15516 20301
rect 16592 18290 16620 20301
rect 17696 18290 17724 20301
rect 7932 18284 7984 18290
rect 7932 18226 7984 18232
rect 9128 18284 9180 18290
rect 9128 18226 9180 18232
rect 9956 18284 10008 18290
rect 9956 18226 10008 18232
rect 11060 18284 11112 18290
rect 11060 18226 11112 18232
rect 11152 18284 11204 18290
rect 11152 18226 11204 18232
rect 12164 18284 12216 18290
rect 12164 18226 12216 18232
rect 13268 18284 13320 18290
rect 13268 18226 13320 18232
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 15476 18284 15528 18290
rect 15476 18226 15528 18232
rect 16580 18284 16632 18290
rect 16580 18226 16632 18232
rect 17684 18284 17736 18290
rect 17684 18226 17736 18232
rect 11072 18170 11100 18226
rect 11980 18216 12032 18222
rect 11072 18142 11192 18170
rect 11980 18158 12032 18164
rect 8484 18080 8536 18086
rect 8484 18022 8536 18028
rect 9956 18080 10008 18086
rect 9956 18022 10008 18028
rect 10048 18080 10100 18086
rect 10048 18022 10100 18028
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 7916 17980 8292 17989
rect 7972 17978 7996 17980
rect 8052 17978 8076 17980
rect 8132 17978 8156 17980
rect 8212 17978 8236 17980
rect 7972 17926 7982 17978
rect 8226 17926 8236 17978
rect 7972 17924 7996 17926
rect 8052 17924 8076 17926
rect 8132 17924 8156 17926
rect 8212 17924 8236 17926
rect 7916 17915 8292 17924
rect 7104 17332 7156 17338
rect 7104 17274 7156 17280
rect 8496 17270 8524 18022
rect 9772 17740 9824 17746
rect 9772 17682 9824 17688
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 8656 17436 9032 17445
rect 8712 17434 8736 17436
rect 8792 17434 8816 17436
rect 8872 17434 8896 17436
rect 8952 17434 8976 17436
rect 8712 17382 8722 17434
rect 8966 17382 8976 17434
rect 8712 17380 8736 17382
rect 8792 17380 8816 17382
rect 8872 17380 8896 17382
rect 8952 17380 8976 17382
rect 8656 17371 9032 17380
rect 9140 17338 9168 17614
rect 9784 17592 9812 17682
rect 9784 17564 9904 17592
rect 9128 17332 9180 17338
rect 9128 17274 9180 17280
rect 8484 17264 8536 17270
rect 8484 17206 8536 17212
rect 7916 16892 8292 16901
rect 7972 16890 7996 16892
rect 8052 16890 8076 16892
rect 8132 16890 8156 16892
rect 8212 16890 8236 16892
rect 7972 16838 7982 16890
rect 8226 16838 8236 16890
rect 7972 16836 7996 16838
rect 8052 16836 8076 16838
rect 8132 16836 8156 16838
rect 8212 16836 8236 16838
rect 7916 16827 8292 16836
rect 9140 16658 9168 17274
rect 9220 17264 9272 17270
rect 9220 17206 9272 17212
rect 9232 16794 9260 17206
rect 9876 17134 9904 17564
rect 9864 17128 9916 17134
rect 9864 17070 9916 17076
rect 9220 16788 9272 16794
rect 9220 16730 9272 16736
rect 9876 16658 9904 17070
rect 9968 16794 9996 18022
rect 10060 17746 10088 18022
rect 10048 17740 10100 17746
rect 10048 17682 10100 17688
rect 11072 17610 11100 18022
rect 11060 17604 11112 17610
rect 11060 17546 11112 17552
rect 11164 17338 11192 18142
rect 11796 18080 11848 18086
rect 11796 18022 11848 18028
rect 11428 17604 11480 17610
rect 11428 17546 11480 17552
rect 11152 17332 11204 17338
rect 11152 17274 11204 17280
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 9128 16652 9180 16658
rect 9128 16594 9180 16600
rect 9864 16652 9916 16658
rect 9864 16594 9916 16600
rect 10140 16652 10192 16658
rect 10140 16594 10192 16600
rect 8656 16348 9032 16357
rect 8712 16346 8736 16348
rect 8792 16346 8816 16348
rect 8872 16346 8896 16348
rect 8952 16346 8976 16348
rect 8712 16294 8722 16346
rect 8966 16294 8976 16346
rect 8712 16292 8736 16294
rect 8792 16292 8816 16294
rect 8872 16292 8896 16294
rect 8952 16292 8976 16294
rect 8656 16283 9032 16292
rect 7288 16244 7340 16250
rect 7288 16186 7340 16192
rect 7840 16244 7892 16250
rect 7840 16186 7892 16192
rect 7300 16114 7328 16186
rect 7104 16108 7156 16114
rect 7288 16108 7340 16114
rect 7156 16068 7288 16096
rect 7104 16050 7156 16056
rect 7288 16050 7340 16056
rect 7748 15972 7800 15978
rect 7748 15914 7800 15920
rect 7012 15632 7064 15638
rect 7012 15574 7064 15580
rect 7024 15434 7052 15574
rect 7472 15564 7524 15570
rect 7472 15506 7524 15512
rect 7012 15428 7064 15434
rect 7012 15370 7064 15376
rect 6920 15360 6972 15366
rect 6920 15302 6972 15308
rect 6932 15094 6960 15302
rect 6920 15088 6972 15094
rect 6920 15030 6972 15036
rect 7024 14890 7052 15370
rect 7484 15026 7512 15506
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7668 15026 7696 15438
rect 7760 15094 7788 15914
rect 7852 15162 7880 16186
rect 9588 16176 9640 16182
rect 9588 16118 9640 16124
rect 8852 16108 8904 16114
rect 8852 16050 8904 16056
rect 7916 15804 8292 15813
rect 7972 15802 7996 15804
rect 8052 15802 8076 15804
rect 8132 15802 8156 15804
rect 8212 15802 8236 15804
rect 7972 15750 7982 15802
rect 8226 15750 8236 15802
rect 7972 15748 7996 15750
rect 8052 15748 8076 15750
rect 8132 15748 8156 15750
rect 8212 15748 8236 15750
rect 7916 15739 8292 15748
rect 8864 15706 8892 16050
rect 9600 15910 9628 16118
rect 9588 15904 9640 15910
rect 9588 15846 9640 15852
rect 8852 15700 8904 15706
rect 8852 15642 8904 15648
rect 9220 15564 9272 15570
rect 9220 15506 9272 15512
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 7840 15156 7892 15162
rect 7840 15098 7892 15104
rect 7748 15088 7800 15094
rect 7748 15030 7800 15036
rect 8312 15026 8340 15302
rect 8656 15260 9032 15269
rect 8712 15258 8736 15260
rect 8792 15258 8816 15260
rect 8872 15258 8896 15260
rect 8952 15258 8976 15260
rect 8712 15206 8722 15258
rect 8966 15206 8976 15258
rect 8712 15204 8736 15206
rect 8792 15204 8816 15206
rect 8872 15204 8896 15206
rect 8952 15204 8976 15206
rect 8656 15195 9032 15204
rect 9140 15094 9168 15438
rect 9232 15366 9260 15506
rect 9600 15502 9628 15846
rect 9588 15496 9640 15502
rect 9588 15438 9640 15444
rect 9956 15496 10008 15502
rect 9956 15438 10008 15444
rect 9220 15360 9272 15366
rect 9220 15302 9272 15308
rect 9128 15088 9180 15094
rect 9128 15030 9180 15036
rect 7472 15020 7524 15026
rect 7472 14962 7524 14968
rect 7656 15020 7708 15026
rect 7656 14962 7708 14968
rect 8300 15020 8352 15026
rect 8300 14962 8352 14968
rect 7012 14884 7064 14890
rect 7012 14826 7064 14832
rect 8668 14816 8720 14822
rect 8668 14758 8720 14764
rect 8760 14816 8812 14822
rect 8760 14758 8812 14764
rect 7916 14716 8292 14725
rect 7972 14714 7996 14716
rect 8052 14714 8076 14716
rect 8132 14714 8156 14716
rect 8212 14714 8236 14716
rect 7972 14662 7982 14714
rect 8226 14662 8236 14714
rect 7972 14660 7996 14662
rect 8052 14660 8076 14662
rect 8132 14660 8156 14662
rect 8212 14660 8236 14662
rect 7916 14651 8292 14660
rect 8680 14618 8708 14758
rect 8668 14612 8720 14618
rect 8668 14554 8720 14560
rect 8772 14414 8800 14758
rect 9232 14618 9260 15302
rect 9600 15162 9628 15438
rect 9588 15156 9640 15162
rect 9588 15098 9640 15104
rect 9968 14958 9996 15438
rect 9956 14952 10008 14958
rect 9956 14894 10008 14900
rect 9220 14612 9272 14618
rect 9220 14554 9272 14560
rect 9864 14476 9916 14482
rect 9864 14418 9916 14424
rect 6828 14408 6880 14414
rect 6828 14350 6880 14356
rect 8760 14408 8812 14414
rect 8760 14350 8812 14356
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 6840 13870 6868 14350
rect 6920 14340 6972 14346
rect 6920 14282 6972 14288
rect 6932 13938 6960 14282
rect 8656 14172 9032 14181
rect 8712 14170 8736 14172
rect 8792 14170 8816 14172
rect 8872 14170 8896 14172
rect 8952 14170 8976 14172
rect 8712 14118 8722 14170
rect 8966 14118 8976 14170
rect 8712 14116 8736 14118
rect 8792 14116 8816 14118
rect 8872 14116 8896 14118
rect 8952 14116 8976 14118
rect 8656 14107 9032 14116
rect 9784 14074 9812 14350
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9876 13938 9904 14418
rect 6920 13932 6972 13938
rect 6920 13874 6972 13880
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9864 13932 9916 13938
rect 9864 13874 9916 13880
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6932 12714 6960 13874
rect 9312 13864 9364 13870
rect 9312 13806 9364 13812
rect 8484 13728 8536 13734
rect 8484 13670 8536 13676
rect 7916 13628 8292 13637
rect 7972 13626 7996 13628
rect 8052 13626 8076 13628
rect 8132 13626 8156 13628
rect 8212 13626 8236 13628
rect 7972 13574 7982 13626
rect 8226 13574 8236 13626
rect 7972 13572 7996 13574
rect 8052 13572 8076 13574
rect 8132 13572 8156 13574
rect 8212 13572 8236 13574
rect 7916 13563 8292 13572
rect 7656 13524 7708 13530
rect 7656 13466 7708 13472
rect 7104 13320 7156 13326
rect 7104 13262 7156 13268
rect 7564 13320 7616 13326
rect 7564 13262 7616 13268
rect 6920 12708 6972 12714
rect 6920 12650 6972 12656
rect 7116 12442 7144 13262
rect 7576 12986 7604 13262
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 7668 12374 7696 13466
rect 7748 13388 7800 13394
rect 7748 13330 7800 13336
rect 7760 12850 7788 13330
rect 8496 12850 8524 13670
rect 8656 13084 9032 13093
rect 8712 13082 8736 13084
rect 8792 13082 8816 13084
rect 8872 13082 8896 13084
rect 8952 13082 8976 13084
rect 8712 13030 8722 13082
rect 8966 13030 8976 13082
rect 8712 13028 8736 13030
rect 8792 13028 8816 13030
rect 8872 13028 8896 13030
rect 8952 13028 8976 13030
rect 8656 13019 9032 13028
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 8484 12844 8536 12850
rect 8484 12786 8536 12792
rect 9324 12782 9352 13806
rect 9508 13394 9536 13874
rect 9588 13796 9640 13802
rect 9588 13738 9640 13744
rect 9496 13388 9548 13394
rect 9496 13330 9548 13336
rect 9508 12782 9536 13330
rect 9600 12986 9628 13738
rect 10152 13326 10180 16594
rect 11164 16522 11192 16934
rect 11152 16516 11204 16522
rect 11152 16458 11204 16464
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10428 15366 10456 15438
rect 11244 15428 11296 15434
rect 11244 15370 11296 15376
rect 10416 15360 10468 15366
rect 10416 15302 10468 15308
rect 10508 15360 10560 15366
rect 10508 15302 10560 15308
rect 10428 15162 10456 15302
rect 10416 15156 10468 15162
rect 10416 15098 10468 15104
rect 10520 15094 10548 15302
rect 10508 15088 10560 15094
rect 10508 15030 10560 15036
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 10876 14952 10928 14958
rect 10876 14894 10928 14900
rect 10888 14618 10916 14894
rect 11060 14816 11112 14822
rect 11060 14758 11112 14764
rect 11072 14618 11100 14758
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 11060 14612 11112 14618
rect 11060 14554 11112 14560
rect 10888 14414 10916 14554
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 10876 14408 10928 14414
rect 10876 14350 10928 14356
rect 10704 13870 10732 14350
rect 11072 14074 11100 14554
rect 11164 14414 11192 14962
rect 11256 14618 11284 15370
rect 11244 14612 11296 14618
rect 11244 14554 11296 14560
rect 11152 14408 11204 14414
rect 11152 14350 11204 14356
rect 10968 14068 11020 14074
rect 10968 14010 11020 14016
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 10980 13954 11008 14010
rect 10980 13926 11100 13954
rect 10692 13864 10744 13870
rect 10692 13806 10744 13812
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 9680 13252 9732 13258
rect 9680 13194 9732 13200
rect 9588 12980 9640 12986
rect 9588 12922 9640 12928
rect 9692 12918 9720 13194
rect 10152 12986 10180 13262
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 9680 12912 9732 12918
rect 9680 12854 9732 12860
rect 9312 12776 9364 12782
rect 9312 12718 9364 12724
rect 9496 12776 9548 12782
rect 9496 12718 9548 12724
rect 7916 12540 8292 12549
rect 7972 12538 7996 12540
rect 8052 12538 8076 12540
rect 8132 12538 8156 12540
rect 8212 12538 8236 12540
rect 7972 12486 7982 12538
rect 8226 12486 8236 12538
rect 7972 12484 7996 12486
rect 8052 12484 8076 12486
rect 8132 12484 8156 12486
rect 8212 12484 8236 12486
rect 7916 12475 8292 12484
rect 7656 12368 7708 12374
rect 7656 12310 7708 12316
rect 7564 12164 7616 12170
rect 7564 12106 7616 12112
rect 6644 12096 6696 12102
rect 6644 12038 6696 12044
rect 7576 11898 7604 12106
rect 8656 11996 9032 12005
rect 8712 11994 8736 11996
rect 8792 11994 8816 11996
rect 8872 11994 8896 11996
rect 8952 11994 8976 11996
rect 8712 11942 8722 11994
rect 8966 11942 8976 11994
rect 8712 11940 8736 11942
rect 8792 11940 8816 11942
rect 8872 11940 8896 11942
rect 8952 11940 8976 11942
rect 8656 11931 9032 11940
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 8484 11756 8536 11762
rect 8484 11698 8536 11704
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 6932 11286 6960 11698
rect 6920 11280 6972 11286
rect 6920 11222 6972 11228
rect 7024 11150 7052 11698
rect 8404 11626 8432 11698
rect 8392 11620 8444 11626
rect 8392 11562 8444 11568
rect 7916 11452 8292 11461
rect 7972 11450 7996 11452
rect 8052 11450 8076 11452
rect 8132 11450 8156 11452
rect 8212 11450 8236 11452
rect 7972 11398 7982 11450
rect 8226 11398 8236 11450
rect 7972 11396 7996 11398
rect 8052 11396 8076 11398
rect 8132 11396 8156 11398
rect 8212 11396 8236 11398
rect 7916 11387 8292 11396
rect 8404 11150 8432 11562
rect 8496 11218 8524 11698
rect 8484 11212 8536 11218
rect 8484 11154 8536 11160
rect 8864 11150 8892 11698
rect 9324 11626 9352 12718
rect 9312 11620 9364 11626
rect 9312 11562 9364 11568
rect 7012 11144 7064 11150
rect 7012 11086 7064 11092
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 8852 11144 8904 11150
rect 8852 11086 8904 11092
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 8484 11076 8536 11082
rect 8484 11018 8536 11024
rect 6644 10736 6696 10742
rect 6644 10678 6696 10684
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 5724 10600 5776 10606
rect 5724 10542 5776 10548
rect 6656 10266 6684 10678
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 3884 10192 3936 10198
rect 3884 10134 3936 10140
rect 3896 9722 3924 10134
rect 4252 9988 4304 9994
rect 4252 9930 4304 9936
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 3976 9580 4028 9586
rect 3976 9522 4028 9528
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 3700 9512 3752 9518
rect 3700 9454 3752 9460
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3988 8974 4016 9522
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 4080 8906 4108 9522
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 4172 9382 4200 9454
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 4264 9178 4292 9930
rect 5724 9648 5776 9654
rect 5724 9590 5776 9596
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 4896 9580 4948 9586
rect 4896 9522 4948 9528
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 4436 9512 4488 9518
rect 4436 9454 4488 9460
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4172 9058 4200 9114
rect 4448 9058 4476 9454
rect 4172 9030 4476 9058
rect 4724 9042 4752 9522
rect 4712 9036 4764 9042
rect 4068 8900 4120 8906
rect 4068 8842 4120 8848
rect 3976 8832 4028 8838
rect 3976 8774 4028 8780
rect 3988 8430 4016 8774
rect 4172 8498 4200 9030
rect 4712 8978 4764 8984
rect 4908 8974 4936 9522
rect 5092 9364 5120 9522
rect 5264 9376 5316 9382
rect 5092 9336 5264 9364
rect 5264 9318 5316 9324
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 5276 8906 5304 9318
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5264 8900 5316 8906
rect 5264 8842 5316 8848
rect 5276 8634 5304 8842
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 3424 8424 3476 8430
rect 3424 8366 3476 8372
rect 3976 8424 4028 8430
rect 3976 8366 4028 8372
rect 3424 7812 3476 7818
rect 3424 7754 3476 7760
rect 3436 7342 3464 7754
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 3792 7268 3844 7274
rect 3792 7210 3844 7216
rect 3804 6798 3832 7210
rect 3896 6798 3924 7346
rect 4172 6866 4200 8434
rect 5184 8294 5212 8434
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5184 7886 5212 8230
rect 5368 7954 5396 8434
rect 5552 8022 5580 8910
rect 5644 8498 5672 8910
rect 5736 8906 5764 9590
rect 6932 9178 6960 11018
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 5724 8900 5776 8906
rect 5724 8842 5776 8848
rect 5736 8634 5764 8842
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5540 8016 5592 8022
rect 5540 7958 5592 7964
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 4160 6860 4212 6866
rect 4160 6802 4212 6808
rect 4724 6798 4752 7142
rect 4816 6934 4844 7346
rect 4804 6928 4856 6934
rect 4804 6870 4856 6876
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 3608 6724 3660 6730
rect 3608 6666 3660 6672
rect 3620 6254 3648 6666
rect 3804 6458 3832 6734
rect 5828 6458 5856 7346
rect 3792 6452 3844 6458
rect 3792 6394 3844 6400
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 6734 6352 6790 6361
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 5908 6316 5960 6322
rect 6734 6287 6736 6296
rect 5908 6258 5960 6264
rect 6788 6287 6790 6296
rect 6736 6258 6788 6264
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 4264 5914 4292 6258
rect 4356 5914 4384 6258
rect 5920 5914 5948 6258
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 5908 5908 5960 5914
rect 5908 5850 5960 5856
rect 6380 5846 6408 6054
rect 7116 5846 7144 10542
rect 7916 10364 8292 10373
rect 7972 10362 7996 10364
rect 8052 10362 8076 10364
rect 8132 10362 8156 10364
rect 8212 10362 8236 10364
rect 7972 10310 7982 10362
rect 8226 10310 8236 10362
rect 7972 10308 7996 10310
rect 8052 10308 8076 10310
rect 8132 10308 8156 10310
rect 8212 10308 8236 10310
rect 7916 10299 8292 10308
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7300 8974 7328 9318
rect 7916 9276 8292 9285
rect 7972 9274 7996 9276
rect 8052 9274 8076 9276
rect 8132 9274 8156 9276
rect 8212 9274 8236 9276
rect 7972 9222 7982 9274
rect 8226 9222 8236 9274
rect 7972 9220 7996 9222
rect 8052 9220 8076 9222
rect 8132 9220 8156 9222
rect 8212 9220 8236 9222
rect 7916 9211 8292 9220
rect 8404 9178 8432 9454
rect 8496 9178 8524 11018
rect 8656 10908 9032 10917
rect 8712 10906 8736 10908
rect 8792 10906 8816 10908
rect 8872 10906 8896 10908
rect 8952 10906 8976 10908
rect 8712 10854 8722 10906
rect 8966 10854 8976 10906
rect 8712 10852 8736 10854
rect 8792 10852 8816 10854
rect 8872 10852 8896 10854
rect 8952 10852 8976 10854
rect 8656 10843 9032 10852
rect 9692 10470 9720 12854
rect 10704 12714 10732 13806
rect 11072 13394 11100 13926
rect 11164 13530 11192 14350
rect 11244 13932 11296 13938
rect 11244 13874 11296 13880
rect 11152 13524 11204 13530
rect 11152 13466 11204 13472
rect 11060 13388 11112 13394
rect 11112 13348 11192 13376
rect 11060 13330 11112 13336
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 10692 12708 10744 12714
rect 10692 12650 10744 12656
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 9680 10464 9732 10470
rect 9680 10406 9732 10412
rect 8656 9820 9032 9829
rect 8712 9818 8736 9820
rect 8792 9818 8816 9820
rect 8872 9818 8896 9820
rect 8952 9818 8976 9820
rect 8712 9766 8722 9818
rect 8966 9766 8976 9818
rect 8712 9764 8736 9766
rect 8792 9764 8816 9766
rect 8872 9764 8896 9766
rect 8952 9764 8976 9766
rect 8656 9755 9032 9764
rect 9692 9654 9720 10406
rect 9784 10198 9812 11698
rect 10520 11218 10548 11698
rect 10796 11354 10824 11698
rect 10784 11348 10836 11354
rect 10784 11290 10836 11296
rect 10508 11212 10560 11218
rect 10508 11154 10560 11160
rect 10692 11008 10744 11014
rect 10692 10950 10744 10956
rect 9772 10192 9824 10198
rect 9772 10134 9824 10140
rect 10704 10130 10732 10950
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 10796 10198 10824 10542
rect 10876 10464 10928 10470
rect 10876 10406 10928 10412
rect 10784 10192 10836 10198
rect 10784 10134 10836 10140
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10048 10056 10100 10062
rect 10048 9998 10100 10004
rect 9772 9988 9824 9994
rect 9772 9930 9824 9936
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 9784 9586 9812 9930
rect 10060 9926 10088 9998
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 10060 9518 10088 9862
rect 10704 9586 10732 10066
rect 10888 10062 10916 10406
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10980 9926 11008 10542
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 10048 9512 10100 9518
rect 10048 9454 10100 9460
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 9496 9376 9548 9382
rect 9496 9318 9548 9324
rect 8392 9172 8444 9178
rect 8392 9114 8444 9120
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8680 8974 8708 9318
rect 9232 9042 9260 9318
rect 9220 9036 9272 9042
rect 9220 8978 9272 8984
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 8668 8968 8720 8974
rect 8668 8910 8720 8916
rect 7380 8900 7432 8906
rect 7380 8842 7432 8848
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 7208 8022 7236 8434
rect 7392 8362 7420 8842
rect 8656 8732 9032 8741
rect 8712 8730 8736 8732
rect 8792 8730 8816 8732
rect 8872 8730 8896 8732
rect 8952 8730 8976 8732
rect 8712 8678 8722 8730
rect 8966 8678 8976 8730
rect 8712 8676 8736 8678
rect 8792 8676 8816 8678
rect 8872 8676 8896 8678
rect 8952 8676 8976 8678
rect 8656 8667 9032 8676
rect 9232 8634 9260 8978
rect 9508 8906 9536 9318
rect 9680 9104 9732 9110
rect 9680 9046 9732 9052
rect 9496 8900 9548 8906
rect 9496 8842 9548 8848
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 9692 8498 9720 9046
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 7380 8356 7432 8362
rect 7380 8298 7432 8304
rect 7484 8090 7512 8434
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7668 8022 7696 8434
rect 7916 8188 8292 8197
rect 7972 8186 7996 8188
rect 8052 8186 8076 8188
rect 8132 8186 8156 8188
rect 8212 8186 8236 8188
rect 7972 8134 7982 8186
rect 8226 8134 8236 8186
rect 7972 8132 7996 8134
rect 8052 8132 8076 8134
rect 8132 8132 8156 8134
rect 8212 8132 8236 8134
rect 7916 8123 8292 8132
rect 7196 8016 7248 8022
rect 7196 7958 7248 7964
rect 7380 8016 7432 8022
rect 7380 7958 7432 7964
rect 7656 8016 7708 8022
rect 7656 7958 7708 7964
rect 7392 7886 7420 7958
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 9496 7880 9548 7886
rect 9496 7822 9548 7828
rect 7852 6905 7880 7822
rect 8656 7644 9032 7653
rect 8712 7642 8736 7644
rect 8792 7642 8816 7644
rect 8872 7642 8896 7644
rect 8952 7642 8976 7644
rect 8712 7590 8722 7642
rect 8966 7590 8976 7642
rect 8712 7588 8736 7590
rect 8792 7588 8816 7590
rect 8872 7588 8896 7590
rect 8952 7588 8976 7590
rect 8656 7579 9032 7588
rect 9508 7546 9536 7822
rect 9600 7546 9628 8434
rect 9692 8022 9720 8434
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 9968 8090 9996 8366
rect 10140 8288 10192 8294
rect 10140 8230 10192 8236
rect 10152 8090 10180 8230
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 9680 8016 9732 8022
rect 9680 7958 9732 7964
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9968 7410 9996 7890
rect 10140 7812 10192 7818
rect 10140 7754 10192 7760
rect 10152 7546 10180 7754
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 9956 7404 10008 7410
rect 9956 7346 10008 7352
rect 7916 7100 8292 7109
rect 7972 7098 7996 7100
rect 8052 7098 8076 7100
rect 8132 7098 8156 7100
rect 8212 7098 8236 7100
rect 7972 7046 7982 7098
rect 8226 7046 8236 7098
rect 7972 7044 7996 7046
rect 8052 7044 8076 7046
rect 8132 7044 8156 7046
rect 8212 7044 8236 7046
rect 7916 7035 8292 7044
rect 7838 6896 7894 6905
rect 9784 6866 9812 7346
rect 9968 7290 9996 7346
rect 9876 7274 9996 7290
rect 9864 7268 9996 7274
rect 9916 7262 9996 7268
rect 9864 7210 9916 7216
rect 9968 7002 9996 7262
rect 9956 6996 10008 7002
rect 9956 6938 10008 6944
rect 10600 6996 10652 7002
rect 10600 6938 10652 6944
rect 7838 6831 7894 6840
rect 9128 6860 9180 6866
rect 9128 6802 9180 6808
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7562 6760 7618 6769
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 6368 5840 6420 5846
rect 6368 5782 6420 5788
rect 7104 5840 7156 5846
rect 7104 5782 7156 5788
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 4172 5234 4200 5510
rect 4448 5302 4476 5646
rect 4436 5296 4488 5302
rect 4436 5238 4488 5244
rect 4632 5234 4660 5646
rect 6644 5636 6696 5642
rect 6644 5578 6696 5584
rect 5816 5364 5868 5370
rect 5816 5306 5868 5312
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 4172 4282 4200 5170
rect 5460 4826 5488 5170
rect 5828 5030 5856 5306
rect 5908 5296 5960 5302
rect 5908 5238 5960 5244
rect 5920 5166 5948 5238
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 4160 4276 4212 4282
rect 4160 4218 4212 4224
rect 3516 4140 3568 4146
rect 3516 4082 3568 4088
rect 3240 3528 3292 3534
rect 3240 3470 3292 3476
rect 2412 3188 2464 3194
rect 2412 3130 2464 3136
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 3148 3188 3200 3194
rect 3148 3130 3200 3136
rect 2884 2990 2912 3130
rect 2872 2984 2924 2990
rect 2872 2926 2924 2932
rect 3252 2854 3280 3470
rect 3424 3120 3476 3126
rect 3424 3062 3476 3068
rect 2320 2848 2372 2854
rect 2320 2790 2372 2796
rect 3240 2848 3292 2854
rect 3240 2790 3292 2796
rect 1916 2748 2292 2757
rect 1972 2746 1996 2748
rect 2052 2746 2076 2748
rect 2132 2746 2156 2748
rect 2212 2746 2236 2748
rect 1972 2694 1982 2746
rect 2226 2694 2236 2746
rect 1972 2692 1996 2694
rect 2052 2692 2076 2694
rect 2132 2692 2156 2694
rect 2212 2692 2236 2694
rect 1916 2683 2292 2692
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 2332 2378 2360 2790
rect 3436 2650 3464 3062
rect 3528 2990 3556 4082
rect 5920 4010 5948 5102
rect 6656 5030 6684 5578
rect 6644 5024 6696 5030
rect 6644 4966 6696 4972
rect 6368 4616 6420 4622
rect 6368 4558 6420 4564
rect 6184 4480 6236 4486
rect 6184 4422 6236 4428
rect 6196 4146 6224 4422
rect 6092 4140 6144 4146
rect 6092 4082 6144 4088
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 4528 4004 4580 4010
rect 4528 3946 4580 3952
rect 5908 4004 5960 4010
rect 5908 3946 5960 3952
rect 4540 3738 4568 3946
rect 4528 3732 4580 3738
rect 4528 3674 4580 3680
rect 6104 3534 6132 4082
rect 6380 4078 6408 4558
rect 7116 4486 7144 5782
rect 7392 5778 7420 6258
rect 7380 5772 7432 5778
rect 7380 5714 7432 5720
rect 7196 5568 7248 5574
rect 7196 5510 7248 5516
rect 7208 5234 7236 5510
rect 7196 5228 7248 5234
rect 7196 5170 7248 5176
rect 7392 5166 7420 5714
rect 7484 5710 7512 6734
rect 7562 6695 7564 6704
rect 7616 6695 7618 6704
rect 9140 6712 9168 6802
rect 9404 6792 9456 6798
rect 9402 6760 9404 6769
rect 9456 6760 9458 6769
rect 9312 6724 9364 6730
rect 7564 6666 7616 6672
rect 9140 6684 9312 6712
rect 7472 5704 7524 5710
rect 7472 5646 7524 5652
rect 7484 5234 7512 5646
rect 7576 5574 7604 6666
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 7656 6384 7708 6390
rect 7656 6326 7708 6332
rect 7668 5914 7696 6326
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 7748 6248 7800 6254
rect 7748 6190 7800 6196
rect 7760 5914 7788 6190
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 7564 5568 7616 5574
rect 7564 5510 7616 5516
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7380 5160 7432 5166
rect 7380 5102 7432 5108
rect 7196 5092 7248 5098
rect 7196 5034 7248 5040
rect 7208 4554 7236 5034
rect 7196 4548 7248 4554
rect 7196 4490 7248 4496
rect 7104 4480 7156 4486
rect 7104 4422 7156 4428
rect 7208 4146 7236 4490
rect 7484 4146 7512 5170
rect 7576 4690 7604 5510
rect 7668 5166 7696 5850
rect 7852 5692 7880 6054
rect 7916 6012 8292 6021
rect 7972 6010 7996 6012
rect 8052 6010 8076 6012
rect 8132 6010 8156 6012
rect 8212 6010 8236 6012
rect 7972 5958 7982 6010
rect 8226 5958 8236 6010
rect 7972 5956 7996 5958
rect 8052 5956 8076 5958
rect 8132 5956 8156 5958
rect 8212 5956 8236 5958
rect 7916 5947 8292 5956
rect 8208 5840 8260 5846
rect 8208 5782 8260 5788
rect 8220 5710 8248 5782
rect 7932 5704 7984 5710
rect 7852 5664 7932 5692
rect 7932 5646 7984 5652
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8300 5704 8352 5710
rect 8404 5692 8432 6258
rect 8588 6254 8616 6598
rect 8656 6556 9032 6565
rect 8712 6554 8736 6556
rect 8792 6554 8816 6556
rect 8872 6554 8896 6556
rect 8952 6554 8976 6556
rect 8712 6502 8722 6554
rect 8966 6502 8976 6554
rect 8712 6500 8736 6502
rect 8792 6500 8816 6502
rect 8872 6500 8896 6502
rect 8952 6500 8976 6502
rect 8656 6491 9032 6500
rect 8576 6248 8628 6254
rect 8576 6190 8628 6196
rect 8352 5664 8432 5692
rect 8300 5646 8352 5652
rect 8128 5574 8156 5646
rect 8116 5568 8168 5574
rect 8116 5510 8168 5516
rect 8312 5370 8340 5646
rect 9140 5642 9168 6684
rect 9402 6695 9458 6704
rect 9312 6666 9364 6672
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9876 5846 9904 6258
rect 10152 6254 10180 6394
rect 10140 6248 10192 6254
rect 10140 6190 10192 6196
rect 9956 6112 10008 6118
rect 9956 6054 10008 6060
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 9968 5914 9996 6054
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 9220 5840 9272 5846
rect 9220 5782 9272 5788
rect 9864 5840 9916 5846
rect 9864 5782 9916 5788
rect 9128 5636 9180 5642
rect 9128 5578 9180 5584
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 7656 5160 7708 5166
rect 7656 5102 7708 5108
rect 7916 4924 8292 4933
rect 7972 4922 7996 4924
rect 8052 4922 8076 4924
rect 8132 4922 8156 4924
rect 8212 4922 8236 4924
rect 7972 4870 7982 4922
rect 8226 4870 8236 4922
rect 7972 4868 7996 4870
rect 8052 4868 8076 4870
rect 8132 4868 8156 4870
rect 8212 4868 8236 4870
rect 7916 4859 8292 4868
rect 8392 4752 8444 4758
rect 8392 4694 8444 4700
rect 7564 4684 7616 4690
rect 7564 4626 7616 4632
rect 7656 4480 7708 4486
rect 7656 4422 7708 4428
rect 6920 4140 6972 4146
rect 7196 4140 7248 4146
rect 6972 4100 7196 4128
rect 6920 4082 6972 4088
rect 7196 4082 7248 4088
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 6368 4072 6420 4078
rect 6368 4014 6420 4020
rect 6552 4004 6604 4010
rect 6552 3946 6604 3952
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 6380 3602 6408 3878
rect 6564 3670 6592 3946
rect 6552 3664 6604 3670
rect 6552 3606 6604 3612
rect 6368 3596 6420 3602
rect 6368 3538 6420 3544
rect 6092 3528 6144 3534
rect 6092 3470 6144 3476
rect 4252 3460 4304 3466
rect 4252 3402 4304 3408
rect 7104 3460 7156 3466
rect 7104 3402 7156 3408
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 3804 2514 3832 3130
rect 3896 3126 3924 3334
rect 3884 3120 3936 3126
rect 3884 3062 3936 3068
rect 4264 2990 4292 3402
rect 5264 3120 5316 3126
rect 5264 3062 5316 3068
rect 3884 2984 3936 2990
rect 3884 2926 3936 2932
rect 4252 2984 4304 2990
rect 4252 2926 4304 2932
rect 3896 2774 3924 2926
rect 3896 2746 4016 2774
rect 3792 2508 3844 2514
rect 3792 2450 3844 2456
rect 3988 2446 4016 2746
rect 5276 2650 5304 3062
rect 7116 3058 7144 3402
rect 7484 3126 7512 4082
rect 7668 4010 7696 4422
rect 8404 4146 8432 4694
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 7656 4004 7708 4010
rect 7656 3946 7708 3952
rect 7668 3534 7696 3946
rect 7916 3836 8292 3845
rect 7972 3834 7996 3836
rect 8052 3834 8076 3836
rect 8132 3834 8156 3836
rect 8212 3834 8236 3836
rect 7972 3782 7982 3834
rect 8226 3782 8236 3834
rect 7972 3780 7996 3782
rect 8052 3780 8076 3782
rect 8132 3780 8156 3782
rect 8212 3780 8236 3782
rect 7916 3771 8292 3780
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8312 3602 8340 3674
rect 8404 3670 8432 4082
rect 8392 3664 8444 3670
rect 8392 3606 8444 3612
rect 8496 3602 8524 5510
rect 8656 5468 9032 5477
rect 8712 5466 8736 5468
rect 8792 5466 8816 5468
rect 8872 5466 8896 5468
rect 8952 5466 8976 5468
rect 8712 5414 8722 5466
rect 8966 5414 8976 5466
rect 8712 5412 8736 5414
rect 8792 5412 8816 5414
rect 8872 5412 8896 5414
rect 8952 5412 8976 5414
rect 8656 5403 9032 5412
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 8680 5030 8708 5306
rect 9140 5234 9168 5578
rect 9232 5370 9260 5782
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9784 5574 9812 5646
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 9220 5364 9272 5370
rect 9220 5306 9272 5312
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 8668 5024 8720 5030
rect 8668 4966 8720 4972
rect 9140 4758 9168 5170
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 9496 5160 9548 5166
rect 9496 5102 9548 5108
rect 9128 4752 9180 4758
rect 9128 4694 9180 4700
rect 9232 4622 9260 5102
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 9324 4690 9352 4966
rect 9312 4684 9364 4690
rect 9312 4626 9364 4632
rect 9508 4622 9536 5102
rect 10060 4826 10088 6054
rect 10152 5234 10180 6190
rect 10416 5908 10468 5914
rect 10416 5850 10468 5856
rect 10232 5840 10284 5846
rect 10232 5782 10284 5788
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 10244 5030 10272 5782
rect 10324 5772 10376 5778
rect 10324 5714 10376 5720
rect 10336 5574 10364 5714
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 10336 5370 10364 5510
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 10428 5234 10456 5850
rect 10612 5846 10640 6938
rect 10690 6216 10746 6225
rect 10690 6151 10746 6160
rect 10600 5840 10652 5846
rect 10600 5782 10652 5788
rect 10704 5642 10732 6151
rect 10692 5636 10744 5642
rect 10692 5578 10744 5584
rect 10876 5568 10928 5574
rect 10876 5510 10928 5516
rect 10416 5228 10468 5234
rect 10416 5170 10468 5176
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 10232 5024 10284 5030
rect 10232 4966 10284 4972
rect 10048 4820 10100 4826
rect 10048 4762 10100 4768
rect 10520 4758 10548 5170
rect 10704 4826 10732 5170
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 10508 4752 10560 4758
rect 10508 4694 10560 4700
rect 8576 4616 8628 4622
rect 8576 4558 8628 4564
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 9496 4616 9548 4622
rect 9496 4558 9548 4564
rect 10692 4616 10744 4622
rect 10796 4604 10824 5170
rect 10888 4690 10916 5510
rect 10980 5098 11008 9862
rect 11072 7954 11100 12922
rect 11164 12918 11192 13348
rect 11152 12912 11204 12918
rect 11152 12854 11204 12860
rect 11152 12776 11204 12782
rect 11152 12718 11204 12724
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 11072 7002 11100 7346
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 11164 5914 11192 12718
rect 11256 12646 11284 13874
rect 11336 13796 11388 13802
rect 11336 13738 11388 13744
rect 11348 13326 11376 13738
rect 11336 13320 11388 13326
rect 11336 13262 11388 13268
rect 11348 12782 11376 13262
rect 11336 12776 11388 12782
rect 11336 12718 11388 12724
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 11336 9580 11388 9586
rect 11336 9522 11388 9528
rect 11348 8498 11376 9522
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 11244 7336 11296 7342
rect 11244 7278 11296 7284
rect 11152 5908 11204 5914
rect 11152 5850 11204 5856
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 10968 5092 11020 5098
rect 10968 5034 11020 5040
rect 10876 4684 10928 4690
rect 10876 4626 10928 4632
rect 10744 4576 10824 4604
rect 10692 4558 10744 4564
rect 8588 4282 8616 4558
rect 8656 4380 9032 4389
rect 8712 4378 8736 4380
rect 8792 4378 8816 4380
rect 8872 4378 8896 4380
rect 8952 4378 8976 4380
rect 8712 4326 8722 4378
rect 8966 4326 8976 4378
rect 8712 4324 8736 4326
rect 8792 4324 8816 4326
rect 8872 4324 8896 4326
rect 8952 4324 8976 4326
rect 8656 4315 9032 4324
rect 8576 4276 8628 4282
rect 8576 4218 8628 4224
rect 9508 4146 9536 4558
rect 9496 4140 9548 4146
rect 9496 4082 9548 4088
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 9770 4040 9826 4049
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 8312 3126 8340 3538
rect 7472 3120 7524 3126
rect 7472 3062 7524 3068
rect 8300 3120 8352 3126
rect 8300 3062 8352 3068
rect 8496 3058 8524 3538
rect 8680 3466 8708 4014
rect 9770 3975 9826 3984
rect 9784 3602 9812 3975
rect 10704 3738 10732 4558
rect 10876 4276 10928 4282
rect 10876 4218 10928 4224
rect 10784 4004 10836 4010
rect 10784 3946 10836 3952
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 8668 3460 8720 3466
rect 8668 3402 8720 3408
rect 8656 3292 9032 3301
rect 8712 3290 8736 3292
rect 8792 3290 8816 3292
rect 8872 3290 8896 3292
rect 8952 3290 8976 3292
rect 8712 3238 8722 3290
rect 8966 3238 8976 3290
rect 8712 3236 8736 3238
rect 8792 3236 8816 3238
rect 8872 3236 8896 3238
rect 8952 3236 8976 3238
rect 8656 3227 9032 3236
rect 9416 3194 9444 3470
rect 9404 3188 9456 3194
rect 9404 3130 9456 3136
rect 9784 3126 9812 3538
rect 10600 3528 10652 3534
rect 10600 3470 10652 3476
rect 10140 3392 10192 3398
rect 10140 3334 10192 3340
rect 9772 3120 9824 3126
rect 9772 3062 9824 3068
rect 10152 3058 10180 3334
rect 10612 3194 10640 3470
rect 10600 3188 10652 3194
rect 10600 3130 10652 3136
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 10140 3052 10192 3058
rect 10140 2994 10192 3000
rect 7564 2916 7616 2922
rect 7564 2858 7616 2864
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 3976 2440 4028 2446
rect 3976 2382 4028 2388
rect 7576 2378 7604 2858
rect 7916 2748 8292 2757
rect 7972 2746 7996 2748
rect 8052 2746 8076 2748
rect 8132 2746 8156 2748
rect 8212 2746 8236 2748
rect 7972 2694 7982 2746
rect 8226 2694 8236 2746
rect 7972 2692 7996 2694
rect 8052 2692 8076 2694
rect 8132 2692 8156 2694
rect 8212 2692 8236 2694
rect 7916 2683 8292 2692
rect 9692 2650 9720 2994
rect 10796 2854 10824 3946
rect 10888 3126 10916 4218
rect 10876 3120 10928 3126
rect 10876 3062 10928 3068
rect 10876 2984 10928 2990
rect 10876 2926 10928 2932
rect 10888 2854 10916 2926
rect 11072 2922 11100 5510
rect 11152 5296 11204 5302
rect 11152 5238 11204 5244
rect 11164 4690 11192 5238
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 11256 4282 11284 7278
rect 11244 4276 11296 4282
rect 11244 4218 11296 4224
rect 11348 4049 11376 8434
rect 11440 7274 11468 17546
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 11716 15706 11744 15846
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 11612 15632 11664 15638
rect 11612 15574 11664 15580
rect 11624 15502 11652 15574
rect 11612 15496 11664 15502
rect 11612 15438 11664 15444
rect 11624 14074 11652 15438
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11612 12912 11664 12918
rect 11612 12854 11664 12860
rect 11624 11830 11652 12854
rect 11612 11824 11664 11830
rect 11612 11766 11664 11772
rect 11624 11626 11652 11766
rect 11612 11620 11664 11626
rect 11612 11562 11664 11568
rect 11624 11150 11652 11562
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11716 11218 11744 11494
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 11624 10674 11652 11086
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11624 9994 11652 10610
rect 11612 9988 11664 9994
rect 11612 9930 11664 9936
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11428 7268 11480 7274
rect 11428 7210 11480 7216
rect 11440 6866 11468 7210
rect 11532 7206 11560 8570
rect 11624 8362 11652 9930
rect 11612 8356 11664 8362
rect 11612 8298 11664 8304
rect 11520 7200 11572 7206
rect 11520 7142 11572 7148
rect 11428 6860 11480 6866
rect 11428 6802 11480 6808
rect 11532 6798 11560 7142
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11532 6186 11560 6734
rect 11612 6724 11664 6730
rect 11612 6666 11664 6672
rect 11624 6322 11652 6666
rect 11612 6316 11664 6322
rect 11612 6258 11664 6264
rect 11520 6180 11572 6186
rect 11520 6122 11572 6128
rect 11716 5370 11744 11154
rect 11808 7954 11836 18022
rect 11992 13394 12020 18158
rect 12164 18148 12216 18154
rect 12164 18090 12216 18096
rect 12176 17610 12204 18090
rect 12440 18080 12492 18086
rect 12438 18048 12440 18057
rect 13268 18080 13320 18086
rect 12492 18048 12494 18057
rect 13268 18022 13320 18028
rect 15476 18080 15528 18086
rect 15476 18022 15528 18028
rect 15568 18080 15620 18086
rect 15568 18022 15620 18028
rect 16028 18080 16080 18086
rect 16028 18022 16080 18028
rect 17224 18080 17276 18086
rect 17224 18022 17276 18028
rect 12438 17983 12494 17992
rect 12164 17604 12216 17610
rect 12164 17546 12216 17552
rect 12624 17604 12676 17610
rect 12624 17546 12676 17552
rect 12256 17536 12308 17542
rect 12256 17478 12308 17484
rect 12348 17536 12400 17542
rect 12348 17478 12400 17484
rect 12072 17128 12124 17134
rect 12072 17070 12124 17076
rect 12084 15609 12112 17070
rect 12268 16114 12296 17478
rect 12360 17202 12388 17478
rect 12636 17338 12664 17546
rect 12624 17332 12676 17338
rect 12624 17274 12676 17280
rect 12348 17196 12400 17202
rect 12348 17138 12400 17144
rect 13280 17134 13308 18022
rect 13916 17980 14292 17989
rect 13972 17978 13996 17980
rect 14052 17978 14076 17980
rect 14132 17978 14156 17980
rect 14212 17978 14236 17980
rect 13972 17926 13982 17978
rect 14226 17926 14236 17978
rect 13972 17924 13996 17926
rect 14052 17924 14076 17926
rect 14132 17924 14156 17926
rect 14212 17924 14236 17926
rect 13916 17915 14292 17924
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 13452 17604 13504 17610
rect 13372 17564 13452 17592
rect 13268 17128 13320 17134
rect 13268 17070 13320 17076
rect 12992 16584 13044 16590
rect 12992 16526 13044 16532
rect 12440 16516 12492 16522
rect 12440 16458 12492 16464
rect 12348 16244 12400 16250
rect 12348 16186 12400 16192
rect 12256 16108 12308 16114
rect 12256 16050 12308 16056
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 12070 15600 12126 15609
rect 12070 15535 12126 15544
rect 12176 15026 12204 15846
rect 12164 15020 12216 15026
rect 12164 14962 12216 14968
rect 12268 14618 12296 16050
rect 12360 15502 12388 16186
rect 12452 15502 12480 16458
rect 12808 16448 12860 16454
rect 12808 16390 12860 16396
rect 12532 16176 12584 16182
rect 12584 16136 12664 16164
rect 12532 16118 12584 16124
rect 12636 15638 12664 16136
rect 12820 16114 12848 16390
rect 13004 16114 13032 16526
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 13372 16046 13400 17564
rect 13452 17546 13504 17552
rect 13556 17270 13584 17682
rect 14556 17672 14608 17678
rect 14556 17614 14608 17620
rect 14280 17536 14332 17542
rect 14280 17478 14332 17484
rect 14292 17270 14320 17478
rect 13544 17264 13596 17270
rect 13544 17206 13596 17212
rect 14280 17264 14332 17270
rect 14280 17206 14332 17212
rect 13556 16658 13584 17206
rect 14568 17202 14596 17614
rect 14656 17436 15032 17445
rect 14712 17434 14736 17436
rect 14792 17434 14816 17436
rect 14872 17434 14896 17436
rect 14952 17434 14976 17436
rect 14712 17382 14722 17434
rect 14966 17382 14976 17434
rect 14712 17380 14736 17382
rect 14792 17380 14816 17382
rect 14872 17380 14896 17382
rect 14952 17380 14976 17382
rect 14656 17371 15032 17380
rect 14556 17196 14608 17202
rect 14556 17138 14608 17144
rect 13916 16892 14292 16901
rect 13972 16890 13996 16892
rect 14052 16890 14076 16892
rect 14132 16890 14156 16892
rect 14212 16890 14236 16892
rect 13972 16838 13982 16890
rect 14226 16838 14236 16890
rect 13972 16836 13996 16838
rect 14052 16836 14076 16838
rect 14132 16836 14156 16838
rect 14212 16836 14236 16838
rect 13916 16827 14292 16836
rect 13912 16720 13964 16726
rect 13912 16662 13964 16668
rect 13544 16652 13596 16658
rect 13544 16594 13596 16600
rect 13452 16448 13504 16454
rect 13452 16390 13504 16396
rect 13084 16040 13136 16046
rect 13084 15982 13136 15988
rect 13360 16040 13412 16046
rect 13360 15982 13412 15988
rect 12624 15632 12676 15638
rect 12624 15574 12676 15580
rect 12714 15600 12770 15609
rect 12636 15502 12664 15574
rect 12714 15535 12770 15544
rect 12728 15502 12756 15535
rect 12348 15496 12400 15502
rect 12348 15438 12400 15444
rect 12440 15496 12492 15502
rect 12440 15438 12492 15444
rect 12624 15496 12676 15502
rect 12624 15438 12676 15444
rect 12716 15496 12768 15502
rect 12768 15456 12848 15484
rect 12716 15438 12768 15444
rect 12256 14612 12308 14618
rect 12256 14554 12308 14560
rect 12360 13920 12388 15438
rect 12452 15008 12480 15438
rect 12532 15360 12584 15366
rect 12532 15302 12584 15308
rect 12544 15162 12572 15302
rect 12532 15156 12584 15162
rect 12532 15098 12584 15104
rect 12452 14980 12572 15008
rect 12360 13892 12480 13920
rect 12348 13796 12400 13802
rect 12268 13756 12348 13784
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 11992 12850 12020 13330
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 12072 13184 12124 13190
rect 12072 13126 12124 13132
rect 11980 12844 12032 12850
rect 11980 12786 12032 12792
rect 12084 12782 12112 13126
rect 12072 12776 12124 12782
rect 12072 12718 12124 12724
rect 11980 9512 12032 9518
rect 11980 9454 12032 9460
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11900 8566 11928 9318
rect 11992 9042 12020 9454
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 12084 9178 12112 9318
rect 12072 9172 12124 9178
rect 12072 9114 12124 9120
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 11888 8560 11940 8566
rect 11888 8502 11940 8508
rect 12072 8424 12124 8430
rect 12072 8366 12124 8372
rect 12084 7954 12112 8366
rect 11796 7948 11848 7954
rect 11796 7890 11848 7896
rect 12072 7948 12124 7954
rect 12072 7890 12124 7896
rect 12084 7342 12112 7890
rect 12176 7410 12204 13262
rect 12268 8566 12296 13756
rect 12348 13738 12400 13744
rect 12452 12986 12480 13892
rect 12544 13802 12572 14980
rect 12532 13796 12584 13802
rect 12532 13738 12584 13744
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12636 12850 12664 15438
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 12728 15026 12756 15302
rect 12820 15026 12848 15456
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12808 15020 12860 15026
rect 12808 14962 12860 14968
rect 12728 13190 12756 14962
rect 12820 14822 12848 14962
rect 13096 14890 13124 15982
rect 13360 15904 13412 15910
rect 13360 15846 13412 15852
rect 13372 15502 13400 15846
rect 13360 15496 13412 15502
rect 13360 15438 13412 15444
rect 13176 15428 13228 15434
rect 13176 15370 13228 15376
rect 13188 15162 13216 15370
rect 13176 15156 13228 15162
rect 13176 15098 13228 15104
rect 13372 14958 13400 15438
rect 13176 14952 13228 14958
rect 13176 14894 13228 14900
rect 13360 14952 13412 14958
rect 13360 14894 13412 14900
rect 13084 14884 13136 14890
rect 13084 14826 13136 14832
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 13084 13932 13136 13938
rect 13084 13874 13136 13880
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12624 12844 12676 12850
rect 12624 12786 12676 12792
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12544 11762 12572 12038
rect 12532 11756 12584 11762
rect 12532 11698 12584 11704
rect 12636 11694 12664 12786
rect 12728 11898 12756 13126
rect 12820 12850 12848 13330
rect 12900 12980 12952 12986
rect 12900 12922 12952 12928
rect 12808 12844 12860 12850
rect 12808 12786 12860 12792
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12820 11778 12848 12786
rect 12728 11762 12848 11778
rect 12912 11762 12940 12922
rect 13096 12850 13124 13874
rect 13188 13410 13216 14894
rect 13360 14612 13412 14618
rect 13360 14554 13412 14560
rect 13268 14068 13320 14074
rect 13268 14010 13320 14016
rect 13280 13530 13308 14010
rect 13372 13938 13400 14554
rect 13464 14074 13492 16390
rect 13556 14414 13584 16594
rect 13924 16590 13952 16662
rect 13912 16584 13964 16590
rect 13912 16526 13964 16532
rect 13924 16114 13952 16526
rect 15108 16448 15160 16454
rect 15108 16390 15160 16396
rect 14656 16348 15032 16357
rect 14712 16346 14736 16348
rect 14792 16346 14816 16348
rect 14872 16346 14896 16348
rect 14952 16346 14976 16348
rect 14712 16294 14722 16346
rect 14966 16294 14976 16346
rect 14712 16292 14736 16294
rect 14792 16292 14816 16294
rect 14872 16292 14896 16294
rect 14952 16292 14976 16294
rect 14656 16283 15032 16292
rect 15120 16250 15148 16390
rect 14004 16244 14056 16250
rect 14004 16186 14056 16192
rect 14464 16244 14516 16250
rect 14464 16186 14516 16192
rect 14832 16244 14884 16250
rect 14832 16186 14884 16192
rect 15108 16244 15160 16250
rect 15108 16186 15160 16192
rect 14016 16114 14044 16186
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 14004 16108 14056 16114
rect 14004 16050 14056 16056
rect 13820 15972 13872 15978
rect 13820 15914 13872 15920
rect 13636 15700 13688 15706
rect 13636 15642 13688 15648
rect 13648 15094 13676 15642
rect 13832 15434 13860 15914
rect 13916 15804 14292 15813
rect 13972 15802 13996 15804
rect 14052 15802 14076 15804
rect 14132 15802 14156 15804
rect 14212 15802 14236 15804
rect 13972 15750 13982 15802
rect 14226 15750 14236 15802
rect 13972 15748 13996 15750
rect 14052 15748 14076 15750
rect 14132 15748 14156 15750
rect 14212 15748 14236 15750
rect 13916 15739 14292 15748
rect 14096 15564 14148 15570
rect 14096 15506 14148 15512
rect 13820 15428 13872 15434
rect 13820 15370 13872 15376
rect 13636 15088 13688 15094
rect 13636 15030 13688 15036
rect 13544 14408 13596 14414
rect 13544 14350 13596 14356
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 13268 13524 13320 13530
rect 13268 13466 13320 13472
rect 13188 13382 13308 13410
rect 13084 12844 13136 12850
rect 13084 12786 13136 12792
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 13084 11892 13136 11898
rect 13084 11834 13136 11840
rect 12716 11756 12848 11762
rect 12768 11750 12848 11756
rect 12900 11756 12952 11762
rect 12716 11698 12768 11704
rect 12900 11698 12952 11704
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 12636 11098 12664 11630
rect 12728 11218 12756 11698
rect 12716 11212 12768 11218
rect 12716 11154 12768 11160
rect 12452 9382 12480 11086
rect 12636 11070 12848 11098
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12728 10062 12756 10202
rect 12532 10056 12584 10062
rect 12716 10056 12768 10062
rect 12584 10016 12664 10044
rect 12532 9998 12584 10004
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12544 9586 12572 9862
rect 12636 9722 12664 10016
rect 12716 9998 12768 10004
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12636 9178 12664 9522
rect 12624 9172 12676 9178
rect 12624 9114 12676 9120
rect 12728 8974 12756 9862
rect 12820 9450 12848 11070
rect 12912 10198 12940 11698
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 13004 11218 13032 11494
rect 12992 11212 13044 11218
rect 12992 11154 13044 11160
rect 12900 10192 12952 10198
rect 12900 10134 12952 10140
rect 13096 10062 13124 11834
rect 13188 11694 13216 12038
rect 13176 11688 13228 11694
rect 13176 11630 13228 11636
rect 13084 10056 13136 10062
rect 13084 9998 13136 10004
rect 12992 9988 13044 9994
rect 12992 9930 13044 9936
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 12912 9586 12940 9862
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 13004 9518 13032 9930
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 13096 9586 13124 9658
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 13188 9518 13216 11630
rect 13280 11150 13308 13382
rect 13372 12918 13400 13874
rect 13464 12986 13492 14010
rect 13556 13326 13584 14350
rect 13544 13320 13596 13326
rect 13544 13262 13596 13268
rect 13544 13184 13596 13190
rect 13544 13126 13596 13132
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 13360 12912 13412 12918
rect 13360 12854 13412 12860
rect 13268 11144 13320 11150
rect 13268 11086 13320 11092
rect 13372 11082 13400 12854
rect 13464 11694 13492 12922
rect 13452 11688 13504 11694
rect 13452 11630 13504 11636
rect 13464 11150 13492 11630
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 13360 11076 13412 11082
rect 13360 11018 13412 11024
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 12992 9512 13044 9518
rect 12992 9454 13044 9460
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 12808 9444 12860 9450
rect 12808 9386 12860 9392
rect 12820 9042 12848 9386
rect 12808 9036 12860 9042
rect 12808 8978 12860 8984
rect 13188 8974 13216 9454
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 13176 8968 13228 8974
rect 13176 8910 13228 8916
rect 13280 8838 13308 10202
rect 13452 10124 13504 10130
rect 13452 10066 13504 10072
rect 13464 9994 13492 10066
rect 13556 10062 13584 13126
rect 13648 12782 13676 15030
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13740 13938 13768 14758
rect 13832 14600 13860 15370
rect 14108 14890 14136 15506
rect 14372 15156 14424 15162
rect 14372 15098 14424 15104
rect 14096 14884 14148 14890
rect 14096 14826 14148 14832
rect 13916 14716 14292 14725
rect 13972 14714 13996 14716
rect 14052 14714 14076 14716
rect 14132 14714 14156 14716
rect 14212 14714 14236 14716
rect 13972 14662 13982 14714
rect 14226 14662 14236 14714
rect 13972 14660 13996 14662
rect 14052 14660 14076 14662
rect 14132 14660 14156 14662
rect 14212 14660 14236 14662
rect 13916 14651 14292 14660
rect 13832 14572 13952 14600
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 13728 13932 13780 13938
rect 13728 13874 13780 13880
rect 13740 13190 13768 13874
rect 13832 13462 13860 14418
rect 13924 13870 13952 14572
rect 14384 14074 14412 15098
rect 14476 15094 14504 16186
rect 14844 16114 14872 16186
rect 14832 16108 14884 16114
rect 14832 16050 14884 16056
rect 14924 16108 14976 16114
rect 14924 16050 14976 16056
rect 14844 15978 14872 16050
rect 14832 15972 14884 15978
rect 14832 15914 14884 15920
rect 14556 15564 14608 15570
rect 14556 15506 14608 15512
rect 14464 15088 14516 15094
rect 14464 15030 14516 15036
rect 14568 15026 14596 15506
rect 14844 15502 14872 15914
rect 14936 15638 14964 16050
rect 15016 16040 15068 16046
rect 15016 15982 15068 15988
rect 15292 16040 15344 16046
rect 15292 15982 15344 15988
rect 14924 15632 14976 15638
rect 14924 15574 14976 15580
rect 14832 15496 14884 15502
rect 14832 15438 14884 15444
rect 14924 15496 14976 15502
rect 15028 15450 15056 15982
rect 15108 15632 15160 15638
rect 15108 15574 15160 15580
rect 15120 15502 15148 15574
rect 14976 15444 15056 15450
rect 14924 15438 15056 15444
rect 15108 15496 15160 15502
rect 15108 15438 15160 15444
rect 14936 15422 15056 15438
rect 14936 15366 14964 15422
rect 14924 15360 14976 15366
rect 14924 15302 14976 15308
rect 14656 15260 15032 15269
rect 14712 15258 14736 15260
rect 14792 15258 14816 15260
rect 14872 15258 14896 15260
rect 14952 15258 14976 15260
rect 14712 15206 14722 15258
rect 14966 15206 14976 15258
rect 14712 15204 14736 15206
rect 14792 15204 14816 15206
rect 14872 15204 14896 15206
rect 14952 15204 14976 15206
rect 14656 15195 15032 15204
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 15120 14958 15148 15438
rect 15304 15162 15332 15982
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 14648 14952 14700 14958
rect 14648 14894 14700 14900
rect 15108 14952 15160 14958
rect 15108 14894 15160 14900
rect 14660 14822 14688 14894
rect 15304 14822 15332 15098
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 14648 14816 14700 14822
rect 14648 14758 14700 14764
rect 15108 14816 15160 14822
rect 15108 14758 15160 14764
rect 15292 14816 15344 14822
rect 15292 14758 15344 14764
rect 14656 14172 15032 14181
rect 14712 14170 14736 14172
rect 14792 14170 14816 14172
rect 14872 14170 14896 14172
rect 14952 14170 14976 14172
rect 14712 14118 14722 14170
rect 14966 14118 14976 14170
rect 14712 14116 14736 14118
rect 14792 14116 14816 14118
rect 14872 14116 14896 14118
rect 14952 14116 14976 14118
rect 14656 14107 15032 14116
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 13912 13864 13964 13870
rect 13912 13806 13964 13812
rect 13916 13628 14292 13637
rect 13972 13626 13996 13628
rect 14052 13626 14076 13628
rect 14132 13626 14156 13628
rect 14212 13626 14236 13628
rect 13972 13574 13982 13626
rect 14226 13574 14236 13626
rect 13972 13572 13996 13574
rect 14052 13572 14076 13574
rect 14132 13572 14156 13574
rect 14212 13572 14236 13574
rect 13916 13563 14292 13572
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 13820 13456 13872 13462
rect 13820 13398 13872 13404
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13636 12776 13688 12782
rect 13636 12718 13688 12724
rect 13648 12434 13676 12718
rect 13924 12646 13952 13466
rect 14280 13252 14332 13258
rect 14280 13194 14332 13200
rect 14292 12986 14320 13194
rect 14280 12980 14332 12986
rect 14280 12922 14332 12928
rect 14278 12880 14334 12889
rect 14384 12850 14412 14010
rect 14648 14000 14700 14006
rect 14648 13942 14700 13948
rect 14464 13796 14516 13802
rect 14464 13738 14516 13744
rect 14476 13326 14504 13738
rect 14660 13462 14688 13942
rect 15120 13938 15148 14758
rect 15292 14000 15344 14006
rect 15292 13942 15344 13948
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 14924 13728 14976 13734
rect 14924 13670 14976 13676
rect 14648 13456 14700 13462
rect 14648 13398 14700 13404
rect 14464 13320 14516 13326
rect 14660 13274 14688 13398
rect 14936 13394 14964 13670
rect 14924 13388 14976 13394
rect 14924 13330 14976 13336
rect 14464 13262 14516 13268
rect 14568 13246 14688 13274
rect 14740 13320 14792 13326
rect 14740 13262 14792 13268
rect 14464 13184 14516 13190
rect 14464 13126 14516 13132
rect 14476 12986 14504 13126
rect 14464 12980 14516 12986
rect 14464 12922 14516 12928
rect 14278 12815 14280 12824
rect 14332 12815 14334 12824
rect 14372 12844 14424 12850
rect 14280 12786 14332 12792
rect 14372 12786 14424 12792
rect 13912 12640 13964 12646
rect 14476 12594 14504 12922
rect 13912 12582 13964 12588
rect 14384 12566 14504 12594
rect 13916 12540 14292 12549
rect 13972 12538 13996 12540
rect 14052 12538 14076 12540
rect 14132 12538 14156 12540
rect 14212 12538 14236 12540
rect 13972 12486 13982 12538
rect 14226 12486 14236 12538
rect 13972 12484 13996 12486
rect 14052 12484 14076 12486
rect 14132 12484 14156 12486
rect 14212 12484 14236 12486
rect 13916 12475 14292 12484
rect 13648 12406 13860 12434
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13648 10198 13676 11494
rect 13728 11076 13780 11082
rect 13728 11018 13780 11024
rect 13636 10192 13688 10198
rect 13636 10134 13688 10140
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13452 9988 13504 9994
rect 13452 9930 13504 9936
rect 13464 9586 13492 9930
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 13372 9110 13400 9386
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 13360 9104 13412 9110
rect 13360 9046 13412 9052
rect 12716 8832 12768 8838
rect 12716 8774 12768 8780
rect 13268 8832 13320 8838
rect 13268 8774 13320 8780
rect 12256 8560 12308 8566
rect 12256 8502 12308 8508
rect 12164 7404 12216 7410
rect 12164 7346 12216 7352
rect 12072 7336 12124 7342
rect 12072 7278 12124 7284
rect 12084 6798 12112 7278
rect 12268 6866 12296 8502
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12452 7886 12480 8230
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 12438 7712 12494 7721
rect 12438 7647 12494 7656
rect 12452 7478 12480 7647
rect 12440 7472 12492 7478
rect 12440 7414 12492 7420
rect 12256 6860 12308 6866
rect 12256 6802 12308 6808
rect 12624 6860 12676 6866
rect 12624 6802 12676 6808
rect 12072 6792 12124 6798
rect 12072 6734 12124 6740
rect 12164 6792 12216 6798
rect 12164 6734 12216 6740
rect 12176 6610 12204 6734
rect 11900 6582 12204 6610
rect 11900 6390 11928 6582
rect 11888 6384 11940 6390
rect 11888 6326 11940 6332
rect 12256 6384 12308 6390
rect 12256 6326 12308 6332
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 11808 5710 11836 6190
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 11900 5778 11928 6054
rect 12164 5840 12216 5846
rect 12164 5782 12216 5788
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 11612 4684 11664 4690
rect 11612 4626 11664 4632
rect 11428 4616 11480 4622
rect 11428 4558 11480 4564
rect 11440 4214 11468 4558
rect 11428 4208 11480 4214
rect 11428 4150 11480 4156
rect 11334 4040 11390 4049
rect 11334 3975 11390 3984
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 11164 3126 11192 3878
rect 11256 3534 11284 3878
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 11348 3398 11376 3975
rect 11440 3534 11468 4150
rect 11624 3534 11652 4626
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 11704 3596 11756 3602
rect 11704 3538 11756 3544
rect 11428 3528 11480 3534
rect 11612 3528 11664 3534
rect 11428 3470 11480 3476
rect 11610 3496 11612 3505
rect 11664 3496 11666 3505
rect 11336 3392 11388 3398
rect 11336 3334 11388 3340
rect 11152 3120 11204 3126
rect 11152 3062 11204 3068
rect 11060 2916 11112 2922
rect 11060 2858 11112 2864
rect 10784 2848 10836 2854
rect 10784 2790 10836 2796
rect 10876 2848 10928 2854
rect 10876 2790 10928 2796
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 11440 2446 11468 3470
rect 11610 3431 11666 3440
rect 11716 3194 11744 3538
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 11992 3058 12020 4218
rect 12176 3602 12204 5782
rect 12268 5642 12296 6326
rect 12636 6322 12664 6802
rect 12624 6316 12676 6322
rect 12624 6258 12676 6264
rect 12440 6248 12492 6254
rect 12440 6190 12492 6196
rect 12452 6066 12480 6190
rect 12636 6118 12664 6258
rect 12624 6112 12676 6118
rect 12360 6038 12480 6066
rect 12544 6072 12624 6100
rect 12360 5642 12388 6038
rect 12256 5636 12308 5642
rect 12256 5578 12308 5584
rect 12348 5636 12400 5642
rect 12348 5578 12400 5584
rect 12268 4826 12296 5578
rect 12256 4820 12308 4826
rect 12256 4762 12308 4768
rect 12360 4282 12388 5578
rect 12544 5166 12572 6072
rect 12624 6054 12676 6060
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 12636 5710 12664 5850
rect 12624 5704 12676 5710
rect 12624 5646 12676 5652
rect 12532 5160 12584 5166
rect 12532 5102 12584 5108
rect 12348 4276 12400 4282
rect 12348 4218 12400 4224
rect 12440 4276 12492 4282
rect 12440 4218 12492 4224
rect 12452 4146 12480 4218
rect 12728 4162 12756 8774
rect 13084 8492 13136 8498
rect 13084 8434 13136 8440
rect 13096 6798 13124 8434
rect 13084 6792 13136 6798
rect 13464 6769 13492 9318
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13556 6866 13584 7346
rect 13636 7336 13688 7342
rect 13636 7278 13688 7284
rect 13544 6860 13596 6866
rect 13544 6802 13596 6808
rect 13084 6734 13136 6740
rect 13450 6760 13506 6769
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 12820 5234 12848 6054
rect 12900 5772 12952 5778
rect 12900 5714 12952 5720
rect 12808 5228 12860 5234
rect 12808 5170 12860 5176
rect 12912 5030 12940 5714
rect 12900 5024 12952 5030
rect 12900 4966 12952 4972
rect 12808 4208 12860 4214
rect 12728 4156 12808 4162
rect 12728 4150 12860 4156
rect 12256 4140 12308 4146
rect 12256 4082 12308 4088
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 12728 4134 12848 4150
rect 12268 3738 12296 4082
rect 12440 4004 12492 4010
rect 12440 3946 12492 3952
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 12164 3596 12216 3602
rect 12164 3538 12216 3544
rect 12452 3534 12480 3946
rect 12728 3670 12756 4134
rect 12912 3942 12940 4966
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12716 3664 12768 3670
rect 12716 3606 12768 3612
rect 12900 3664 12952 3670
rect 12900 3606 12952 3612
rect 12912 3534 12940 3606
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 12716 3528 12768 3534
rect 12716 3470 12768 3476
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 12348 3460 12400 3466
rect 12348 3402 12400 3408
rect 12360 3194 12388 3402
rect 12348 3188 12400 3194
rect 12348 3130 12400 3136
rect 12452 3058 12480 3470
rect 12728 3126 12756 3470
rect 12716 3120 12768 3126
rect 12716 3062 12768 3068
rect 11980 3052 12032 3058
rect 11980 2994 12032 3000
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 11992 2922 12020 2994
rect 11980 2916 12032 2922
rect 11980 2858 12032 2864
rect 12728 2854 12756 3062
rect 12912 2990 12940 3470
rect 12900 2984 12952 2990
rect 12900 2926 12952 2932
rect 12348 2848 12400 2854
rect 12348 2790 12400 2796
rect 12716 2848 12768 2854
rect 12716 2790 12768 2796
rect 12360 2446 12388 2790
rect 12728 2446 12756 2790
rect 12912 2582 12940 2926
rect 13096 2774 13124 6734
rect 13450 6695 13506 6704
rect 13464 5778 13492 6695
rect 13452 5772 13504 5778
rect 13452 5714 13504 5720
rect 13452 5636 13504 5642
rect 13452 5578 13504 5584
rect 13360 4548 13412 4554
rect 13360 4490 13412 4496
rect 13176 3732 13228 3738
rect 13176 3674 13228 3680
rect 13004 2746 13124 2774
rect 12900 2576 12952 2582
rect 12900 2518 12952 2524
rect 13004 2514 13032 2746
rect 13188 2650 13216 3674
rect 13372 3398 13400 4490
rect 13464 4282 13492 5578
rect 13452 4276 13504 4282
rect 13452 4218 13504 4224
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 13556 3670 13584 4082
rect 13648 4078 13676 7278
rect 13740 5778 13768 11018
rect 13832 9586 13860 12406
rect 13916 11452 14292 11461
rect 13972 11450 13996 11452
rect 14052 11450 14076 11452
rect 14132 11450 14156 11452
rect 14212 11450 14236 11452
rect 13972 11398 13982 11450
rect 14226 11398 14236 11450
rect 13972 11396 13996 11398
rect 14052 11396 14076 11398
rect 14132 11396 14156 11398
rect 14212 11396 14236 11398
rect 13916 11387 14292 11396
rect 14384 11218 14412 12566
rect 14464 12300 14516 12306
rect 14464 12242 14516 12248
rect 14372 11212 14424 11218
rect 14372 11154 14424 11160
rect 13916 10364 14292 10373
rect 13972 10362 13996 10364
rect 14052 10362 14076 10364
rect 14132 10362 14156 10364
rect 14212 10362 14236 10364
rect 13972 10310 13982 10362
rect 14226 10310 14236 10362
rect 13972 10308 13996 10310
rect 14052 10308 14076 10310
rect 14132 10308 14156 10310
rect 14212 10308 14236 10310
rect 13916 10299 14292 10308
rect 14096 10192 14148 10198
rect 14096 10134 14148 10140
rect 14278 10160 14334 10169
rect 13912 10056 13964 10062
rect 13912 9998 13964 10004
rect 13820 9580 13872 9586
rect 13820 9522 13872 9528
rect 13924 9364 13952 9998
rect 13832 9336 13952 9364
rect 14004 9376 14056 9382
rect 13832 6984 13860 9336
rect 14108 9364 14136 10134
rect 14278 10095 14334 10104
rect 14188 9648 14240 9654
rect 14186 9616 14188 9625
rect 14240 9616 14242 9625
rect 14186 9551 14242 9560
rect 14292 9489 14320 10095
rect 14278 9480 14334 9489
rect 14278 9415 14334 9424
rect 14056 9336 14136 9364
rect 14384 9364 14412 11154
rect 14476 10305 14504 12242
rect 14568 11762 14596 13246
rect 14752 13190 14780 13262
rect 14740 13184 14792 13190
rect 14740 13126 14792 13132
rect 14656 13084 15032 13093
rect 14712 13082 14736 13084
rect 14792 13082 14816 13084
rect 14872 13082 14896 13084
rect 14952 13082 14976 13084
rect 14712 13030 14722 13082
rect 14966 13030 14976 13082
rect 14712 13028 14736 13030
rect 14792 13028 14816 13030
rect 14872 13028 14896 13030
rect 14952 13028 14976 13030
rect 14656 13019 15032 13028
rect 14656 11996 15032 12005
rect 14712 11994 14736 11996
rect 14792 11994 14816 11996
rect 14872 11994 14896 11996
rect 14952 11994 14976 11996
rect 14712 11942 14722 11994
rect 14966 11942 14976 11994
rect 14712 11940 14736 11942
rect 14792 11940 14816 11942
rect 14872 11940 14896 11942
rect 14952 11940 14976 11942
rect 14656 11931 15032 11940
rect 15304 11830 15332 13942
rect 15396 13938 15424 14962
rect 15488 14346 15516 18022
rect 15580 17746 15608 18022
rect 15568 17740 15620 17746
rect 15568 17682 15620 17688
rect 15660 17604 15712 17610
rect 15660 17546 15712 17552
rect 15672 17338 15700 17546
rect 15660 17332 15712 17338
rect 15660 17274 15712 17280
rect 16040 16658 16068 18022
rect 16764 17672 16816 17678
rect 16764 17614 16816 17620
rect 16488 17604 16540 17610
rect 16488 17546 16540 17552
rect 16028 16652 16080 16658
rect 16028 16594 16080 16600
rect 15568 16584 15620 16590
rect 15568 16526 15620 16532
rect 15580 16454 15608 16526
rect 15568 16448 15620 16454
rect 15568 16390 15620 16396
rect 15844 16448 15896 16454
rect 15844 16390 15896 16396
rect 15580 16182 15608 16390
rect 15568 16176 15620 16182
rect 15568 16118 15620 16124
rect 15856 16114 15884 16390
rect 16500 16182 16528 17546
rect 16776 17202 16804 17614
rect 17040 17536 17092 17542
rect 17040 17478 17092 17484
rect 16764 17196 16816 17202
rect 16764 17138 16816 17144
rect 16488 16176 16540 16182
rect 16488 16118 16540 16124
rect 15844 16108 15896 16114
rect 15844 16050 15896 16056
rect 15660 15428 15712 15434
rect 15660 15370 15712 15376
rect 15672 15026 15700 15370
rect 16500 15178 16528 16118
rect 16776 16114 16804 17138
rect 16856 17128 16908 17134
rect 16856 17070 16908 17076
rect 16764 16108 16816 16114
rect 16764 16050 16816 16056
rect 16500 15150 16620 15178
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 16026 14920 16082 14929
rect 15936 14884 15988 14890
rect 16026 14855 16082 14864
rect 15936 14826 15988 14832
rect 15476 14340 15528 14346
rect 15476 14282 15528 14288
rect 15752 14068 15804 14074
rect 15752 14010 15804 14016
rect 15384 13932 15436 13938
rect 15384 13874 15436 13880
rect 15660 13796 15712 13802
rect 15660 13738 15712 13744
rect 15384 13728 15436 13734
rect 15384 13670 15436 13676
rect 15476 13728 15528 13734
rect 15476 13670 15528 13676
rect 15396 13326 15424 13670
rect 15384 13320 15436 13326
rect 15384 13262 15436 13268
rect 15488 12918 15516 13670
rect 15476 12912 15528 12918
rect 15476 12854 15528 12860
rect 15566 12880 15622 12889
rect 15566 12815 15568 12824
rect 15620 12815 15622 12824
rect 15568 12786 15620 12792
rect 15580 12442 15608 12786
rect 15672 12782 15700 13738
rect 15764 12850 15792 14010
rect 15752 12844 15804 12850
rect 15752 12786 15804 12792
rect 15660 12776 15712 12782
rect 15660 12718 15712 12724
rect 15844 12708 15896 12714
rect 15844 12650 15896 12656
rect 15568 12436 15620 12442
rect 15568 12378 15620 12384
rect 15752 12436 15804 12442
rect 15752 12378 15804 12384
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 15292 11824 15344 11830
rect 15292 11766 15344 11772
rect 14556 11756 14608 11762
rect 14556 11698 14608 11704
rect 14462 10296 14518 10305
rect 14462 10231 14518 10240
rect 14464 10192 14516 10198
rect 14464 10134 14516 10140
rect 14476 9518 14504 10134
rect 14568 10062 14596 11698
rect 15108 11688 15160 11694
rect 15108 11630 15160 11636
rect 14656 10908 15032 10917
rect 14712 10906 14736 10908
rect 14792 10906 14816 10908
rect 14872 10906 14896 10908
rect 14952 10906 14976 10908
rect 14712 10854 14722 10906
rect 14966 10854 14976 10906
rect 14712 10852 14736 10854
rect 14792 10852 14816 10854
rect 14872 10852 14896 10854
rect 14952 10852 14976 10854
rect 14656 10843 15032 10852
rect 15120 10810 15148 11630
rect 15304 11150 15332 11766
rect 15672 11762 15700 12038
rect 15764 11762 15792 12378
rect 15856 11898 15884 12650
rect 15844 11892 15896 11898
rect 15844 11834 15896 11840
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 15672 11642 15700 11698
rect 15580 11614 15700 11642
rect 15384 11212 15436 11218
rect 15384 11154 15436 11160
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 15108 10804 15160 10810
rect 15108 10746 15160 10752
rect 14556 10056 14608 10062
rect 14556 9998 14608 10004
rect 14556 9920 14608 9926
rect 14556 9862 14608 9868
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14568 9382 14596 9862
rect 14656 9820 15032 9829
rect 14712 9818 14736 9820
rect 14792 9818 14816 9820
rect 14872 9818 14896 9820
rect 14952 9818 14976 9820
rect 14712 9766 14722 9818
rect 14966 9766 14976 9818
rect 14712 9764 14736 9766
rect 14792 9764 14816 9766
rect 14872 9764 14896 9766
rect 14952 9764 14976 9766
rect 14656 9755 15032 9764
rect 15120 9602 15148 10746
rect 15200 10600 15252 10606
rect 15200 10542 15252 10548
rect 15304 10554 15332 11086
rect 15396 10690 15424 11154
rect 15396 10662 15516 10690
rect 15212 10266 15240 10542
rect 15304 10526 15424 10554
rect 15200 10260 15252 10266
rect 15200 10202 15252 10208
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 14936 9586 15148 9602
rect 15200 9648 15252 9654
rect 15200 9590 15252 9596
rect 14924 9580 15148 9586
rect 14976 9574 15148 9580
rect 14924 9522 14976 9528
rect 15108 9512 15160 9518
rect 15108 9454 15160 9460
rect 14924 9444 14976 9450
rect 14924 9386 14976 9392
rect 14556 9376 14608 9382
rect 14384 9336 14504 9364
rect 14004 9318 14056 9324
rect 13916 9276 14292 9285
rect 13972 9274 13996 9276
rect 14052 9274 14076 9276
rect 14132 9274 14156 9276
rect 14212 9274 14236 9276
rect 13972 9222 13982 9274
rect 14226 9222 14236 9274
rect 13972 9220 13996 9222
rect 14052 9220 14076 9222
rect 14132 9220 14156 9222
rect 14212 9220 14236 9222
rect 13916 9211 14292 9220
rect 14476 9042 14504 9336
rect 14556 9318 14608 9324
rect 14568 9178 14596 9318
rect 14936 9178 14964 9386
rect 15016 9376 15068 9382
rect 15016 9318 15068 9324
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14924 9172 14976 9178
rect 14924 9114 14976 9120
rect 14464 9036 14516 9042
rect 14464 8978 14516 8984
rect 14568 8906 14596 9114
rect 15028 8974 15056 9318
rect 15120 8974 15148 9454
rect 15212 9110 15240 9590
rect 15304 9518 15332 9998
rect 15396 9592 15424 10526
rect 15488 9722 15516 10662
rect 15580 10062 15608 11614
rect 15660 11552 15712 11558
rect 15660 11494 15712 11500
rect 15672 11354 15700 11494
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 15672 10606 15700 11290
rect 15764 11150 15792 11698
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15752 10668 15804 10674
rect 15752 10610 15804 10616
rect 15660 10600 15712 10606
rect 15660 10542 15712 10548
rect 15672 10062 15700 10542
rect 15764 10130 15792 10610
rect 15752 10124 15804 10130
rect 15752 10066 15804 10072
rect 15568 10056 15620 10062
rect 15568 9998 15620 10004
rect 15660 10056 15712 10062
rect 15660 9998 15712 10004
rect 15568 9920 15620 9926
rect 15568 9862 15620 9868
rect 15476 9716 15528 9722
rect 15476 9658 15528 9664
rect 15384 9586 15436 9592
rect 15488 9586 15516 9658
rect 15580 9586 15608 9862
rect 15750 9616 15806 9625
rect 15384 9528 15436 9534
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15568 9580 15620 9586
rect 15568 9522 15620 9528
rect 15660 9580 15712 9586
rect 15750 9551 15752 9560
rect 15660 9522 15712 9528
rect 15804 9551 15806 9560
rect 15752 9522 15804 9528
rect 15292 9512 15344 9518
rect 15292 9454 15344 9460
rect 15304 9110 15332 9454
rect 15200 9104 15252 9110
rect 15200 9046 15252 9052
rect 15292 9104 15344 9110
rect 15292 9046 15344 9052
rect 15212 8974 15240 9046
rect 15016 8968 15068 8974
rect 15016 8910 15068 8916
rect 15108 8968 15160 8974
rect 15108 8910 15160 8916
rect 15200 8968 15252 8974
rect 15200 8910 15252 8916
rect 14556 8900 14608 8906
rect 14556 8842 14608 8848
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 14656 8732 15032 8741
rect 14712 8730 14736 8732
rect 14792 8730 14816 8732
rect 14872 8730 14896 8732
rect 14952 8730 14976 8732
rect 14712 8678 14722 8730
rect 14966 8678 14976 8730
rect 14712 8676 14736 8678
rect 14792 8676 14816 8678
rect 14872 8676 14896 8678
rect 14952 8676 14976 8678
rect 14656 8667 15032 8676
rect 13916 8188 14292 8197
rect 13972 8186 13996 8188
rect 14052 8186 14076 8188
rect 14132 8186 14156 8188
rect 14212 8186 14236 8188
rect 13972 8134 13982 8186
rect 14226 8134 14236 8186
rect 13972 8132 13996 8134
rect 14052 8132 14076 8134
rect 14132 8132 14156 8134
rect 14212 8132 14236 8134
rect 13916 8123 14292 8132
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 14372 7812 14424 7818
rect 14372 7754 14424 7760
rect 14384 7410 14412 7754
rect 14372 7404 14424 7410
rect 14372 7346 14424 7352
rect 13916 7100 14292 7109
rect 13972 7098 13996 7100
rect 14052 7098 14076 7100
rect 14132 7098 14156 7100
rect 14212 7098 14236 7100
rect 13972 7046 13982 7098
rect 14226 7046 14236 7098
rect 13972 7044 13996 7046
rect 14052 7044 14076 7046
rect 14132 7044 14156 7046
rect 14212 7044 14236 7046
rect 13916 7035 14292 7044
rect 14384 7002 14412 7346
rect 14476 7342 14504 7822
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 14372 6996 14424 7002
rect 13832 6956 13952 6984
rect 13820 6792 13872 6798
rect 13820 6734 13872 6740
rect 13728 5772 13780 5778
rect 13728 5714 13780 5720
rect 13740 5370 13768 5714
rect 13832 5370 13860 6734
rect 13924 6662 13952 6956
rect 14372 6938 14424 6944
rect 14370 6896 14426 6905
rect 14370 6831 14372 6840
rect 14424 6831 14426 6840
rect 14372 6802 14424 6808
rect 14568 6798 14596 7686
rect 14656 7644 15032 7653
rect 14712 7642 14736 7644
rect 14792 7642 14816 7644
rect 14872 7642 14896 7644
rect 14952 7642 14976 7644
rect 14712 7590 14722 7642
rect 14966 7590 14976 7642
rect 14712 7588 14736 7590
rect 14792 7588 14816 7590
rect 14872 7588 14896 7590
rect 14952 7588 14976 7590
rect 14656 7579 15032 7588
rect 15120 7478 15148 8774
rect 15108 7472 15160 7478
rect 15108 7414 15160 7420
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 14004 6792 14056 6798
rect 14002 6760 14004 6769
rect 14556 6792 14608 6798
rect 14056 6760 14058 6769
rect 14556 6734 14608 6740
rect 14660 6730 14688 7278
rect 14740 6792 14792 6798
rect 14740 6734 14792 6740
rect 15016 6792 15068 6798
rect 15120 6780 15148 7414
rect 15200 6996 15252 7002
rect 15200 6938 15252 6944
rect 15212 6798 15240 6938
rect 15068 6752 15148 6780
rect 15200 6792 15252 6798
rect 15016 6734 15068 6740
rect 15200 6734 15252 6740
rect 15566 6760 15622 6769
rect 14002 6695 14058 6704
rect 14648 6724 14700 6730
rect 14648 6666 14700 6672
rect 14752 6662 14780 6734
rect 15566 6695 15622 6704
rect 13912 6656 13964 6662
rect 13912 6598 13964 6604
rect 14372 6656 14424 6662
rect 14372 6598 14424 6604
rect 14740 6656 14792 6662
rect 14740 6598 14792 6604
rect 15108 6656 15160 6662
rect 15108 6598 15160 6604
rect 14384 6390 14412 6598
rect 14656 6556 15032 6565
rect 14712 6554 14736 6556
rect 14792 6554 14816 6556
rect 14872 6554 14896 6556
rect 14952 6554 14976 6556
rect 14712 6502 14722 6554
rect 14966 6502 14976 6554
rect 14712 6500 14736 6502
rect 14792 6500 14816 6502
rect 14872 6500 14896 6502
rect 14952 6500 14976 6502
rect 14462 6488 14518 6497
rect 14656 6491 15032 6500
rect 14462 6423 14518 6432
rect 14280 6384 14332 6390
rect 14280 6326 14332 6332
rect 14372 6384 14424 6390
rect 14372 6326 14424 6332
rect 14292 6236 14320 6326
rect 14476 6304 14504 6423
rect 14556 6316 14608 6322
rect 14476 6276 14556 6304
rect 14476 6236 14504 6276
rect 14556 6258 14608 6264
rect 14832 6316 14884 6322
rect 14832 6258 14884 6264
rect 14292 6208 14504 6236
rect 14372 6112 14424 6118
rect 14372 6054 14424 6060
rect 13916 6012 14292 6021
rect 13972 6010 13996 6012
rect 14052 6010 14076 6012
rect 14132 6010 14156 6012
rect 14212 6010 14236 6012
rect 13972 5958 13982 6010
rect 14226 5958 14236 6010
rect 13972 5956 13996 5958
rect 14052 5956 14076 5958
rect 14132 5956 14156 5958
rect 14212 5956 14236 5958
rect 13916 5947 14292 5956
rect 14280 5840 14332 5846
rect 14280 5782 14332 5788
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 13740 5166 13768 5306
rect 13728 5160 13780 5166
rect 13728 5102 13780 5108
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 13740 4026 13768 5102
rect 13832 4486 13860 5306
rect 14108 5302 14136 5510
rect 14096 5296 14148 5302
rect 14096 5238 14148 5244
rect 14292 5234 14320 5782
rect 14384 5234 14412 6054
rect 14280 5228 14332 5234
rect 14280 5170 14332 5176
rect 14372 5228 14424 5234
rect 14372 5170 14424 5176
rect 13916 4924 14292 4933
rect 13972 4922 13996 4924
rect 14052 4922 14076 4924
rect 14132 4922 14156 4924
rect 14212 4922 14236 4924
rect 13972 4870 13982 4922
rect 14226 4870 14236 4922
rect 13972 4868 13996 4870
rect 14052 4868 14076 4870
rect 14132 4868 14156 4870
rect 14212 4868 14236 4870
rect 13916 4859 14292 4868
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 14476 4214 14504 6208
rect 14844 5778 14872 6258
rect 14648 5772 14700 5778
rect 14568 5732 14648 5760
rect 14568 5234 14596 5732
rect 14648 5714 14700 5720
rect 14832 5772 14884 5778
rect 14832 5714 14884 5720
rect 14656 5468 15032 5477
rect 14712 5466 14736 5468
rect 14792 5466 14816 5468
rect 14872 5466 14896 5468
rect 14952 5466 14976 5468
rect 14712 5414 14722 5466
rect 14966 5414 14976 5466
rect 14712 5412 14736 5414
rect 14792 5412 14816 5414
rect 14872 5412 14896 5414
rect 14952 5412 14976 5414
rect 14656 5403 15032 5412
rect 14556 5228 14608 5234
rect 14556 5170 14608 5176
rect 14556 5024 14608 5030
rect 14556 4966 14608 4972
rect 14464 4208 14516 4214
rect 14464 4150 14516 4156
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 13544 3664 13596 3670
rect 13544 3606 13596 3612
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 13556 3126 13584 3606
rect 13544 3120 13596 3126
rect 13544 3062 13596 3068
rect 13648 3040 13676 4014
rect 13740 3998 13860 4026
rect 13728 3936 13780 3942
rect 13728 3878 13780 3884
rect 13740 3738 13768 3878
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13832 3534 13860 3998
rect 13916 3836 14292 3845
rect 13972 3834 13996 3836
rect 14052 3834 14076 3836
rect 14132 3834 14156 3836
rect 14212 3834 14236 3836
rect 13972 3782 13982 3834
rect 14226 3782 14236 3834
rect 13972 3780 13996 3782
rect 14052 3780 14076 3782
rect 14132 3780 14156 3782
rect 14212 3780 14236 3782
rect 13916 3771 14292 3780
rect 14384 3738 14412 4082
rect 14568 3942 14596 4966
rect 14656 4380 15032 4389
rect 14712 4378 14736 4380
rect 14792 4378 14816 4380
rect 14872 4378 14896 4380
rect 14952 4378 14976 4380
rect 14712 4326 14722 4378
rect 14966 4326 14976 4378
rect 14712 4324 14736 4326
rect 14792 4324 14816 4326
rect 14872 4324 14896 4326
rect 14952 4324 14976 4326
rect 14656 4315 15032 4324
rect 14832 4276 14884 4282
rect 14832 4218 14884 4224
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14568 3738 14596 3878
rect 14844 3738 14872 4218
rect 15120 4010 15148 6598
rect 15580 5778 15608 6695
rect 15568 5772 15620 5778
rect 15568 5714 15620 5720
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 15292 5228 15344 5234
rect 15292 5170 15344 5176
rect 15304 4078 15332 5170
rect 15396 4078 15424 5646
rect 15568 4684 15620 4690
rect 15568 4626 15620 4632
rect 15292 4072 15344 4078
rect 15292 4014 15344 4020
rect 15384 4072 15436 4078
rect 15384 4014 15436 4020
rect 15108 4004 15160 4010
rect 15108 3946 15160 3952
rect 15476 3936 15528 3942
rect 15476 3878 15528 3884
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 14556 3732 14608 3738
rect 14556 3674 14608 3680
rect 14832 3732 14884 3738
rect 14832 3674 14884 3680
rect 14372 3596 14424 3602
rect 14372 3538 14424 3544
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 13728 3052 13780 3058
rect 13648 3012 13728 3040
rect 13648 2854 13676 3012
rect 13728 2994 13780 3000
rect 14384 2922 14412 3538
rect 15488 3534 15516 3878
rect 15580 3738 15608 4626
rect 15568 3732 15620 3738
rect 15568 3674 15620 3680
rect 15672 3602 15700 9522
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 15752 7880 15804 7886
rect 15752 7822 15804 7828
rect 15764 7546 15792 7822
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15856 7426 15884 8910
rect 15948 7886 15976 14826
rect 16040 14822 16068 14855
rect 16028 14816 16080 14822
rect 16028 14758 16080 14764
rect 16028 13932 16080 13938
rect 16028 13874 16080 13880
rect 16040 11762 16068 13874
rect 16592 13870 16620 15150
rect 16776 15026 16804 16050
rect 16764 15020 16816 15026
rect 16764 14962 16816 14968
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 16684 14346 16712 14758
rect 16672 14340 16724 14346
rect 16672 14282 16724 14288
rect 16868 13938 16896 17070
rect 17052 16522 17080 17478
rect 17040 16516 17092 16522
rect 17040 16458 17092 16464
rect 16948 15904 17000 15910
rect 16948 15846 17000 15852
rect 16960 15434 16988 15846
rect 17236 15570 17264 18022
rect 17224 15564 17276 15570
rect 17224 15506 17276 15512
rect 17500 15496 17552 15502
rect 17500 15438 17552 15444
rect 16948 15428 17000 15434
rect 16948 15370 17000 15376
rect 17512 14482 17540 15438
rect 17500 14476 17552 14482
rect 17500 14418 17552 14424
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 16856 13932 16908 13938
rect 16856 13874 16908 13880
rect 16580 13864 16632 13870
rect 16580 13806 16632 13812
rect 16396 13388 16448 13394
rect 16396 13330 16448 13336
rect 16212 13184 16264 13190
rect 16212 13126 16264 13132
rect 16224 12986 16252 13126
rect 16212 12980 16264 12986
rect 16212 12922 16264 12928
rect 16408 12850 16436 13330
rect 16592 13326 16620 13806
rect 16868 13326 16896 13874
rect 17420 13734 17448 14214
rect 17408 13728 17460 13734
rect 17408 13670 17460 13676
rect 17420 13394 17448 13670
rect 17408 13388 17460 13394
rect 17408 13330 17460 13336
rect 16580 13320 16632 13326
rect 16580 13262 16632 13268
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16856 13320 16908 13326
rect 16856 13262 16908 13268
rect 16120 12844 16172 12850
rect 16120 12786 16172 12792
rect 16396 12844 16448 12850
rect 16396 12786 16448 12792
rect 16132 12102 16160 12786
rect 16592 12782 16620 13262
rect 16776 12850 16804 13262
rect 16764 12844 16816 12850
rect 16868 12832 16896 13262
rect 16948 12844 17000 12850
rect 16868 12804 16948 12832
rect 16764 12786 16816 12792
rect 16948 12786 17000 12792
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 16224 12434 16252 12582
rect 16224 12406 16344 12434
rect 16212 12300 16264 12306
rect 16212 12242 16264 12248
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 16224 11762 16252 12242
rect 16028 11756 16080 11762
rect 16028 11698 16080 11704
rect 16212 11756 16264 11762
rect 16212 11698 16264 11704
rect 16120 11280 16172 11286
rect 16120 11222 16172 11228
rect 16132 11082 16160 11222
rect 16316 11082 16344 12406
rect 16592 11830 16620 12718
rect 16776 12238 16804 12786
rect 16960 12306 16988 12786
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16580 11824 16632 11830
rect 16580 11766 16632 11772
rect 16776 11762 16804 12174
rect 16960 11898 16988 12242
rect 16948 11892 17000 11898
rect 16948 11834 17000 11840
rect 16764 11756 16816 11762
rect 16764 11698 16816 11704
rect 16948 11756 17000 11762
rect 16948 11698 17000 11704
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 16120 11076 16172 11082
rect 16120 11018 16172 11024
rect 16304 11076 16356 11082
rect 16304 11018 16356 11024
rect 16132 9654 16160 11018
rect 16120 9648 16172 9654
rect 16120 9590 16172 9596
rect 16132 9382 16160 9590
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 15936 7880 15988 7886
rect 15936 7822 15988 7828
rect 16212 7744 16264 7750
rect 16212 7686 16264 7692
rect 15764 7398 15884 7426
rect 15764 4146 15792 7398
rect 16224 6798 16252 7686
rect 16212 6792 16264 6798
rect 16212 6734 16264 6740
rect 15936 6180 15988 6186
rect 15936 6122 15988 6128
rect 15948 5302 15976 6122
rect 16224 5914 16252 6734
rect 16316 6458 16344 11018
rect 16580 10736 16632 10742
rect 16580 10678 16632 10684
rect 16592 10441 16620 10678
rect 16776 10674 16804 11086
rect 16672 10668 16724 10674
rect 16672 10610 16724 10616
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 16578 10432 16634 10441
rect 16578 10367 16634 10376
rect 16684 10282 16712 10610
rect 16960 10606 16988 11698
rect 17040 11552 17092 11558
rect 17040 11494 17092 11500
rect 17052 11218 17080 11494
rect 17040 11212 17092 11218
rect 17040 11154 17092 11160
rect 16948 10600 17000 10606
rect 16868 10548 16948 10554
rect 16868 10542 17000 10548
rect 16868 10526 16988 10542
rect 17052 10538 17080 11154
rect 17040 10532 17092 10538
rect 16592 10254 16804 10282
rect 16868 10266 16896 10526
rect 17040 10474 17092 10480
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 16592 10198 16620 10254
rect 16580 10192 16632 10198
rect 16580 10134 16632 10140
rect 16672 10192 16724 10198
rect 16672 10134 16724 10140
rect 16580 9920 16632 9926
rect 16580 9862 16632 9868
rect 16592 9586 16620 9862
rect 16580 9580 16632 9586
rect 16580 9522 16632 9528
rect 16396 8832 16448 8838
rect 16396 8774 16448 8780
rect 16304 6452 16356 6458
rect 16304 6394 16356 6400
rect 16212 5908 16264 5914
rect 16212 5850 16264 5856
rect 16408 5778 16436 8774
rect 16488 7744 16540 7750
rect 16488 7686 16540 7692
rect 16500 7410 16528 7686
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 16486 6352 16542 6361
rect 16486 6287 16542 6296
rect 16500 5914 16528 6287
rect 16684 6225 16712 10134
rect 16776 8906 16804 10254
rect 16856 10260 16908 10266
rect 16856 10202 16908 10208
rect 16960 10062 16988 10406
rect 17052 10062 17080 10474
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 17040 10056 17092 10062
rect 17040 9998 17092 10004
rect 17132 10056 17184 10062
rect 17132 9998 17184 10004
rect 16856 9580 16908 9586
rect 16856 9522 16908 9528
rect 16868 8974 16896 9522
rect 17144 9518 17172 9998
rect 17224 9580 17276 9586
rect 17224 9522 17276 9528
rect 17132 9512 17184 9518
rect 17132 9454 17184 9460
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 17052 9042 17080 9318
rect 17040 9036 17092 9042
rect 17040 8978 17092 8984
rect 17144 8974 17172 9454
rect 17236 9110 17264 9522
rect 17224 9104 17276 9110
rect 17224 9046 17276 9052
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 16764 8900 16816 8906
rect 16764 8842 16816 8848
rect 17144 8634 17172 8910
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 17224 7200 17276 7206
rect 17224 7142 17276 7148
rect 17236 6866 17264 7142
rect 17224 6860 17276 6866
rect 17224 6802 17276 6808
rect 16670 6216 16726 6225
rect 16670 6151 16726 6160
rect 16488 5908 16540 5914
rect 16488 5850 16540 5856
rect 16580 5840 16632 5846
rect 16580 5782 16632 5788
rect 16396 5772 16448 5778
rect 16396 5714 16448 5720
rect 16304 5636 16356 5642
rect 16304 5578 16356 5584
rect 16316 5370 16344 5578
rect 16304 5364 16356 5370
rect 16304 5306 16356 5312
rect 15936 5296 15988 5302
rect 15936 5238 15988 5244
rect 15948 5030 15976 5238
rect 16028 5228 16080 5234
rect 16028 5170 16080 5176
rect 15936 5024 15988 5030
rect 15936 4966 15988 4972
rect 16040 4690 16068 5170
rect 16592 4826 16620 5782
rect 16672 5772 16724 5778
rect 16672 5714 16724 5720
rect 16580 4820 16632 4826
rect 16580 4762 16632 4768
rect 16684 4758 16712 5714
rect 16764 5024 16816 5030
rect 16764 4966 16816 4972
rect 16672 4752 16724 4758
rect 16672 4694 16724 4700
rect 16028 4684 16080 4690
rect 16028 4626 16080 4632
rect 16776 4622 16804 4966
rect 16764 4616 16816 4622
rect 16764 4558 16816 4564
rect 15844 4208 15896 4214
rect 15844 4150 15896 4156
rect 15752 4140 15804 4146
rect 15752 4082 15804 4088
rect 15660 3596 15712 3602
rect 15580 3556 15660 3584
rect 14648 3528 14700 3534
rect 14568 3488 14648 3516
rect 14568 3194 14596 3488
rect 14648 3470 14700 3476
rect 15476 3528 15528 3534
rect 15476 3470 15528 3476
rect 15108 3392 15160 3398
rect 15108 3334 15160 3340
rect 14656 3292 15032 3301
rect 14712 3290 14736 3292
rect 14792 3290 14816 3292
rect 14872 3290 14896 3292
rect 14952 3290 14976 3292
rect 14712 3238 14722 3290
rect 14966 3238 14976 3290
rect 14712 3236 14736 3238
rect 14792 3236 14816 3238
rect 14872 3236 14896 3238
rect 14952 3236 14976 3238
rect 14656 3227 15032 3236
rect 15120 3194 15148 3334
rect 14556 3188 14608 3194
rect 14556 3130 14608 3136
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 15580 3058 15608 3556
rect 15660 3538 15712 3544
rect 15764 3505 15792 4082
rect 15856 3534 15884 4150
rect 15844 3528 15896 3534
rect 15750 3496 15806 3505
rect 15660 3460 15712 3466
rect 15844 3470 15896 3476
rect 15750 3431 15806 3440
rect 15660 3402 15712 3408
rect 15568 3052 15620 3058
rect 15568 2994 15620 3000
rect 15672 2922 15700 3402
rect 15764 3126 15792 3431
rect 15752 3120 15804 3126
rect 15752 3062 15804 3068
rect 14372 2916 14424 2922
rect 14372 2858 14424 2864
rect 15660 2916 15712 2922
rect 15660 2858 15712 2864
rect 13636 2848 13688 2854
rect 13636 2790 13688 2796
rect 13916 2748 14292 2757
rect 13972 2746 13996 2748
rect 14052 2746 14076 2748
rect 14132 2746 14156 2748
rect 14212 2746 14236 2748
rect 13972 2694 13982 2746
rect 14226 2694 14236 2746
rect 13972 2692 13996 2694
rect 14052 2692 14076 2694
rect 14132 2692 14156 2694
rect 14212 2692 14236 2694
rect 13916 2683 14292 2692
rect 13176 2644 13228 2650
rect 13176 2586 13228 2592
rect 12992 2508 13044 2514
rect 12992 2450 13044 2456
rect 9404 2440 9456 2446
rect 9404 2382 9456 2388
rect 11428 2440 11480 2446
rect 11428 2382 11480 2388
rect 12348 2440 12400 2446
rect 12348 2382 12400 2388
rect 12716 2440 12768 2446
rect 12716 2382 12768 2388
rect 2320 2372 2372 2378
rect 2320 2314 2372 2320
rect 7564 2372 7616 2378
rect 7564 2314 7616 2320
rect 1398 2272 1454 2281
rect 1398 2207 1454 2216
rect 2656 2204 3032 2213
rect 2712 2202 2736 2204
rect 2792 2202 2816 2204
rect 2872 2202 2896 2204
rect 2952 2202 2976 2204
rect 2712 2150 2722 2202
rect 2966 2150 2976 2202
rect 2712 2148 2736 2150
rect 2792 2148 2816 2150
rect 2872 2148 2896 2150
rect 2952 2148 2976 2150
rect 2656 2139 3032 2148
rect 8656 2204 9032 2213
rect 8712 2202 8736 2204
rect 8792 2202 8816 2204
rect 8872 2202 8896 2204
rect 8952 2202 8976 2204
rect 8712 2150 8722 2202
rect 8966 2150 8976 2202
rect 8712 2148 8736 2150
rect 8792 2148 8816 2150
rect 8872 2148 8896 2150
rect 8952 2148 8976 2150
rect 8656 2139 9032 2148
rect 9416 800 9444 2382
rect 14656 2204 15032 2213
rect 14712 2202 14736 2204
rect 14792 2202 14816 2204
rect 14872 2202 14896 2204
rect 14952 2202 14976 2204
rect 14712 2150 14722 2202
rect 14966 2150 14976 2202
rect 14712 2148 14736 2150
rect 14792 2148 14816 2150
rect 14872 2148 14896 2150
rect 14952 2148 14976 2150
rect 14656 2139 15032 2148
rect 9402 0 9458 800
<< via2 >>
rect 1214 18536 1270 18592
rect 2656 18522 2712 18524
rect 2736 18522 2792 18524
rect 2816 18522 2872 18524
rect 2896 18522 2952 18524
rect 2976 18522 3032 18524
rect 2656 18470 2658 18522
rect 2658 18470 2710 18522
rect 2710 18470 2712 18522
rect 2736 18470 2774 18522
rect 2774 18470 2786 18522
rect 2786 18470 2792 18522
rect 2816 18470 2838 18522
rect 2838 18470 2850 18522
rect 2850 18470 2872 18522
rect 2896 18470 2902 18522
rect 2902 18470 2914 18522
rect 2914 18470 2952 18522
rect 2976 18470 2978 18522
rect 2978 18470 3030 18522
rect 3030 18470 3032 18522
rect 2656 18468 2712 18470
rect 2736 18468 2792 18470
rect 2816 18468 2872 18470
rect 2896 18468 2952 18470
rect 2976 18468 3032 18470
rect 1916 17978 1972 17980
rect 1996 17978 2052 17980
rect 2076 17978 2132 17980
rect 2156 17978 2212 17980
rect 2236 17978 2292 17980
rect 1916 17926 1918 17978
rect 1918 17926 1970 17978
rect 1970 17926 1972 17978
rect 1996 17926 2034 17978
rect 2034 17926 2046 17978
rect 2046 17926 2052 17978
rect 2076 17926 2098 17978
rect 2098 17926 2110 17978
rect 2110 17926 2132 17978
rect 2156 17926 2162 17978
rect 2162 17926 2174 17978
rect 2174 17926 2212 17978
rect 2236 17926 2238 17978
rect 2238 17926 2290 17978
rect 2290 17926 2292 17978
rect 1916 17924 1972 17926
rect 1996 17924 2052 17926
rect 2076 17924 2132 17926
rect 2156 17924 2212 17926
rect 2236 17924 2292 17926
rect 1306 17448 1362 17504
rect 2656 17434 2712 17436
rect 2736 17434 2792 17436
rect 2816 17434 2872 17436
rect 2896 17434 2952 17436
rect 2976 17434 3032 17436
rect 2656 17382 2658 17434
rect 2658 17382 2710 17434
rect 2710 17382 2712 17434
rect 2736 17382 2774 17434
rect 2774 17382 2786 17434
rect 2786 17382 2792 17434
rect 2816 17382 2838 17434
rect 2838 17382 2850 17434
rect 2850 17382 2872 17434
rect 2896 17382 2902 17434
rect 2902 17382 2914 17434
rect 2914 17382 2952 17434
rect 2976 17382 2978 17434
rect 2978 17382 3030 17434
rect 3030 17382 3032 17434
rect 2656 17380 2712 17382
rect 2736 17380 2792 17382
rect 2816 17380 2872 17382
rect 2896 17380 2952 17382
rect 2976 17380 3032 17382
rect 1916 16890 1972 16892
rect 1996 16890 2052 16892
rect 2076 16890 2132 16892
rect 2156 16890 2212 16892
rect 2236 16890 2292 16892
rect 1916 16838 1918 16890
rect 1918 16838 1970 16890
rect 1970 16838 1972 16890
rect 1996 16838 2034 16890
rect 2034 16838 2046 16890
rect 2046 16838 2052 16890
rect 2076 16838 2098 16890
rect 2098 16838 2110 16890
rect 2110 16838 2132 16890
rect 2156 16838 2162 16890
rect 2162 16838 2174 16890
rect 2174 16838 2212 16890
rect 2236 16838 2238 16890
rect 2238 16838 2290 16890
rect 2290 16838 2292 16890
rect 1916 16836 1972 16838
rect 1996 16836 2052 16838
rect 2076 16836 2132 16838
rect 2156 16836 2212 16838
rect 2236 16836 2292 16838
rect 846 16496 902 16552
rect 2656 16346 2712 16348
rect 2736 16346 2792 16348
rect 2816 16346 2872 16348
rect 2896 16346 2952 16348
rect 2976 16346 3032 16348
rect 2656 16294 2658 16346
rect 2658 16294 2710 16346
rect 2710 16294 2712 16346
rect 2736 16294 2774 16346
rect 2774 16294 2786 16346
rect 2786 16294 2792 16346
rect 2816 16294 2838 16346
rect 2838 16294 2850 16346
rect 2850 16294 2872 16346
rect 2896 16294 2902 16346
rect 2902 16294 2914 16346
rect 2914 16294 2952 16346
rect 2976 16294 2978 16346
rect 2978 16294 3030 16346
rect 3030 16294 3032 16346
rect 2656 16292 2712 16294
rect 2736 16292 2792 16294
rect 2816 16292 2872 16294
rect 2896 16292 2952 16294
rect 2976 16292 3032 16294
rect 846 15408 902 15464
rect 1916 15802 1972 15804
rect 1996 15802 2052 15804
rect 2076 15802 2132 15804
rect 2156 15802 2212 15804
rect 2236 15802 2292 15804
rect 1916 15750 1918 15802
rect 1918 15750 1970 15802
rect 1970 15750 1972 15802
rect 1996 15750 2034 15802
rect 2034 15750 2046 15802
rect 2046 15750 2052 15802
rect 2076 15750 2098 15802
rect 2098 15750 2110 15802
rect 2110 15750 2132 15802
rect 2156 15750 2162 15802
rect 2162 15750 2174 15802
rect 2174 15750 2212 15802
rect 2236 15750 2238 15802
rect 2238 15750 2290 15802
rect 2290 15750 2292 15802
rect 1916 15748 1972 15750
rect 1996 15748 2052 15750
rect 2076 15748 2132 15750
rect 2156 15748 2212 15750
rect 2236 15748 2292 15750
rect 1916 14714 1972 14716
rect 1996 14714 2052 14716
rect 2076 14714 2132 14716
rect 2156 14714 2212 14716
rect 2236 14714 2292 14716
rect 1916 14662 1918 14714
rect 1918 14662 1970 14714
rect 1970 14662 1972 14714
rect 1996 14662 2034 14714
rect 2034 14662 2046 14714
rect 2046 14662 2052 14714
rect 2076 14662 2098 14714
rect 2098 14662 2110 14714
rect 2110 14662 2132 14714
rect 2156 14662 2162 14714
rect 2162 14662 2174 14714
rect 2174 14662 2212 14714
rect 2236 14662 2238 14714
rect 2238 14662 2290 14714
rect 2290 14662 2292 14714
rect 1916 14660 1972 14662
rect 1996 14660 2052 14662
rect 2076 14660 2132 14662
rect 2156 14660 2212 14662
rect 2236 14660 2292 14662
rect 2656 15258 2712 15260
rect 2736 15258 2792 15260
rect 2816 15258 2872 15260
rect 2896 15258 2952 15260
rect 2976 15258 3032 15260
rect 2656 15206 2658 15258
rect 2658 15206 2710 15258
rect 2710 15206 2712 15258
rect 2736 15206 2774 15258
rect 2774 15206 2786 15258
rect 2786 15206 2792 15258
rect 2816 15206 2838 15258
rect 2838 15206 2850 15258
rect 2850 15206 2872 15258
rect 2896 15206 2902 15258
rect 2902 15206 2914 15258
rect 2914 15206 2952 15258
rect 2976 15206 2978 15258
rect 2978 15206 3030 15258
rect 3030 15206 3032 15258
rect 2656 15204 2712 15206
rect 2736 15204 2792 15206
rect 2816 15204 2872 15206
rect 2896 15204 2952 15206
rect 2976 15204 3032 15206
rect 846 14320 902 14376
rect 1916 13626 1972 13628
rect 1996 13626 2052 13628
rect 2076 13626 2132 13628
rect 2156 13626 2212 13628
rect 2236 13626 2292 13628
rect 1916 13574 1918 13626
rect 1918 13574 1970 13626
rect 1970 13574 1972 13626
rect 1996 13574 2034 13626
rect 2034 13574 2046 13626
rect 2046 13574 2052 13626
rect 2076 13574 2098 13626
rect 2098 13574 2110 13626
rect 2110 13574 2132 13626
rect 2156 13574 2162 13626
rect 2162 13574 2174 13626
rect 2174 13574 2212 13626
rect 2236 13574 2238 13626
rect 2238 13574 2290 13626
rect 2290 13574 2292 13626
rect 1916 13572 1972 13574
rect 1996 13572 2052 13574
rect 2076 13572 2132 13574
rect 2156 13572 2212 13574
rect 2236 13572 2292 13574
rect 2656 14170 2712 14172
rect 2736 14170 2792 14172
rect 2816 14170 2872 14172
rect 2896 14170 2952 14172
rect 2976 14170 3032 14172
rect 2656 14118 2658 14170
rect 2658 14118 2710 14170
rect 2710 14118 2712 14170
rect 2736 14118 2774 14170
rect 2774 14118 2786 14170
rect 2786 14118 2792 14170
rect 2816 14118 2838 14170
rect 2838 14118 2850 14170
rect 2850 14118 2872 14170
rect 2896 14118 2902 14170
rect 2902 14118 2914 14170
rect 2914 14118 2952 14170
rect 2976 14118 2978 14170
rect 2978 14118 3030 14170
rect 3030 14118 3032 14170
rect 2656 14116 2712 14118
rect 2736 14116 2792 14118
rect 2816 14116 2872 14118
rect 2896 14116 2952 14118
rect 2976 14116 3032 14118
rect 3238 14864 3294 14920
rect 846 13232 902 13288
rect 1916 12538 1972 12540
rect 1996 12538 2052 12540
rect 2076 12538 2132 12540
rect 2156 12538 2212 12540
rect 2236 12538 2292 12540
rect 1916 12486 1918 12538
rect 1918 12486 1970 12538
rect 1970 12486 1972 12538
rect 1996 12486 2034 12538
rect 2034 12486 2046 12538
rect 2046 12486 2052 12538
rect 2076 12486 2098 12538
rect 2098 12486 2110 12538
rect 2110 12486 2132 12538
rect 2156 12486 2162 12538
rect 2162 12486 2174 12538
rect 2174 12486 2212 12538
rect 2236 12486 2238 12538
rect 2238 12486 2290 12538
rect 2290 12486 2292 12538
rect 1916 12484 1972 12486
rect 1996 12484 2052 12486
rect 2076 12484 2132 12486
rect 2156 12484 2212 12486
rect 2236 12484 2292 12486
rect 2656 13082 2712 13084
rect 2736 13082 2792 13084
rect 2816 13082 2872 13084
rect 2896 13082 2952 13084
rect 2976 13082 3032 13084
rect 2656 13030 2658 13082
rect 2658 13030 2710 13082
rect 2710 13030 2712 13082
rect 2736 13030 2774 13082
rect 2774 13030 2786 13082
rect 2786 13030 2792 13082
rect 2816 13030 2838 13082
rect 2838 13030 2850 13082
rect 2850 13030 2872 13082
rect 2896 13030 2902 13082
rect 2902 13030 2914 13082
rect 2914 13030 2952 13082
rect 2976 13030 2978 13082
rect 2978 13030 3030 13082
rect 3030 13030 3032 13082
rect 2656 13028 2712 13030
rect 2736 13028 2792 13030
rect 2816 13028 2872 13030
rect 2896 13028 2952 13030
rect 2976 13028 3032 13030
rect 846 12144 902 12200
rect 1916 11450 1972 11452
rect 1996 11450 2052 11452
rect 2076 11450 2132 11452
rect 2156 11450 2212 11452
rect 2236 11450 2292 11452
rect 1916 11398 1918 11450
rect 1918 11398 1970 11450
rect 1970 11398 1972 11450
rect 1996 11398 2034 11450
rect 2034 11398 2046 11450
rect 2046 11398 2052 11450
rect 2076 11398 2098 11450
rect 2098 11398 2110 11450
rect 2110 11398 2132 11450
rect 2156 11398 2162 11450
rect 2162 11398 2174 11450
rect 2174 11398 2212 11450
rect 2236 11398 2238 11450
rect 2238 11398 2290 11450
rect 2290 11398 2292 11450
rect 1916 11396 1972 11398
rect 1996 11396 2052 11398
rect 2076 11396 2132 11398
rect 2156 11396 2212 11398
rect 2236 11396 2292 11398
rect 2656 11994 2712 11996
rect 2736 11994 2792 11996
rect 2816 11994 2872 11996
rect 2896 11994 2952 11996
rect 2976 11994 3032 11996
rect 2656 11942 2658 11994
rect 2658 11942 2710 11994
rect 2710 11942 2712 11994
rect 2736 11942 2774 11994
rect 2774 11942 2786 11994
rect 2786 11942 2792 11994
rect 2816 11942 2838 11994
rect 2838 11942 2850 11994
rect 2850 11942 2872 11994
rect 2896 11942 2902 11994
rect 2902 11942 2914 11994
rect 2914 11942 2952 11994
rect 2976 11942 2978 11994
rect 2978 11942 3030 11994
rect 3030 11942 3032 11994
rect 2656 11940 2712 11942
rect 2736 11940 2792 11942
rect 2816 11940 2872 11942
rect 2896 11940 2952 11942
rect 2976 11940 3032 11942
rect 1306 10920 1362 10976
rect 1916 10362 1972 10364
rect 1996 10362 2052 10364
rect 2076 10362 2132 10364
rect 2156 10362 2212 10364
rect 2236 10362 2292 10364
rect 1916 10310 1918 10362
rect 1918 10310 1970 10362
rect 1970 10310 1972 10362
rect 1996 10310 2034 10362
rect 2034 10310 2046 10362
rect 2046 10310 2052 10362
rect 2076 10310 2098 10362
rect 2098 10310 2110 10362
rect 2110 10310 2132 10362
rect 2156 10310 2162 10362
rect 2162 10310 2174 10362
rect 2174 10310 2212 10362
rect 2236 10310 2238 10362
rect 2238 10310 2290 10362
rect 2290 10310 2292 10362
rect 1916 10308 1972 10310
rect 1996 10308 2052 10310
rect 2076 10308 2132 10310
rect 2156 10308 2212 10310
rect 2236 10308 2292 10310
rect 1306 9832 1362 9888
rect 2656 10906 2712 10908
rect 2736 10906 2792 10908
rect 2816 10906 2872 10908
rect 2896 10906 2952 10908
rect 2976 10906 3032 10908
rect 2656 10854 2658 10906
rect 2658 10854 2710 10906
rect 2710 10854 2712 10906
rect 2736 10854 2774 10906
rect 2774 10854 2786 10906
rect 2786 10854 2792 10906
rect 2816 10854 2838 10906
rect 2838 10854 2850 10906
rect 2850 10854 2872 10906
rect 2896 10854 2902 10906
rect 2902 10854 2914 10906
rect 2914 10854 2952 10906
rect 2976 10854 2978 10906
rect 2978 10854 3030 10906
rect 3030 10854 3032 10906
rect 2656 10852 2712 10854
rect 2736 10852 2792 10854
rect 2816 10852 2872 10854
rect 2896 10852 2952 10854
rect 2976 10852 3032 10854
rect 2656 9818 2712 9820
rect 2736 9818 2792 9820
rect 2816 9818 2872 9820
rect 2896 9818 2952 9820
rect 2976 9818 3032 9820
rect 2656 9766 2658 9818
rect 2658 9766 2710 9818
rect 2710 9766 2712 9818
rect 2736 9766 2774 9818
rect 2774 9766 2786 9818
rect 2786 9766 2792 9818
rect 2816 9766 2838 9818
rect 2838 9766 2850 9818
rect 2850 9766 2872 9818
rect 2896 9766 2902 9818
rect 2902 9766 2914 9818
rect 2914 9766 2952 9818
rect 2976 9766 2978 9818
rect 2978 9766 3030 9818
rect 3030 9766 3032 9818
rect 2656 9764 2712 9766
rect 2736 9764 2792 9766
rect 2816 9764 2872 9766
rect 2896 9764 2952 9766
rect 2976 9764 3032 9766
rect 1916 9274 1972 9276
rect 1996 9274 2052 9276
rect 2076 9274 2132 9276
rect 2156 9274 2212 9276
rect 2236 9274 2292 9276
rect 1916 9222 1918 9274
rect 1918 9222 1970 9274
rect 1970 9222 1972 9274
rect 1996 9222 2034 9274
rect 2034 9222 2046 9274
rect 2046 9222 2052 9274
rect 2076 9222 2098 9274
rect 2098 9222 2110 9274
rect 2110 9222 2132 9274
rect 2156 9222 2162 9274
rect 2162 9222 2174 9274
rect 2174 9222 2212 9274
rect 2236 9222 2238 9274
rect 2238 9222 2290 9274
rect 2290 9222 2292 9274
rect 1916 9220 1972 9222
rect 1996 9220 2052 9222
rect 2076 9220 2132 9222
rect 2156 9220 2212 9222
rect 2236 9220 2292 9222
rect 1306 8744 1362 8800
rect 2656 8730 2712 8732
rect 2736 8730 2792 8732
rect 2816 8730 2872 8732
rect 2896 8730 2952 8732
rect 2976 8730 3032 8732
rect 2656 8678 2658 8730
rect 2658 8678 2710 8730
rect 2710 8678 2712 8730
rect 2736 8678 2774 8730
rect 2774 8678 2786 8730
rect 2786 8678 2792 8730
rect 2816 8678 2838 8730
rect 2838 8678 2850 8730
rect 2850 8678 2872 8730
rect 2896 8678 2902 8730
rect 2902 8678 2914 8730
rect 2914 8678 2952 8730
rect 2976 8678 2978 8730
rect 2978 8678 3030 8730
rect 3030 8678 3032 8730
rect 2656 8676 2712 8678
rect 2736 8676 2792 8678
rect 2816 8676 2872 8678
rect 2896 8676 2952 8678
rect 2976 8676 3032 8678
rect 1916 8186 1972 8188
rect 1996 8186 2052 8188
rect 2076 8186 2132 8188
rect 2156 8186 2212 8188
rect 2236 8186 2292 8188
rect 1916 8134 1918 8186
rect 1918 8134 1970 8186
rect 1970 8134 1972 8186
rect 1996 8134 2034 8186
rect 2034 8134 2046 8186
rect 2046 8134 2052 8186
rect 2076 8134 2098 8186
rect 2098 8134 2110 8186
rect 2110 8134 2132 8186
rect 2156 8134 2162 8186
rect 2162 8134 2174 8186
rect 2174 8134 2212 8186
rect 2236 8134 2238 8186
rect 2238 8134 2290 8186
rect 2290 8134 2292 8186
rect 1916 8132 1972 8134
rect 1996 8132 2052 8134
rect 2076 8132 2132 8134
rect 2156 8132 2212 8134
rect 2236 8132 2292 8134
rect 1306 7656 1362 7712
rect 2656 7642 2712 7644
rect 2736 7642 2792 7644
rect 2816 7642 2872 7644
rect 2896 7642 2952 7644
rect 2976 7642 3032 7644
rect 2656 7590 2658 7642
rect 2658 7590 2710 7642
rect 2710 7590 2712 7642
rect 2736 7590 2774 7642
rect 2774 7590 2786 7642
rect 2786 7590 2792 7642
rect 2816 7590 2838 7642
rect 2838 7590 2850 7642
rect 2850 7590 2872 7642
rect 2896 7590 2902 7642
rect 2902 7590 2914 7642
rect 2914 7590 2952 7642
rect 2976 7590 2978 7642
rect 2978 7590 3030 7642
rect 3030 7590 3032 7642
rect 2656 7588 2712 7590
rect 2736 7588 2792 7590
rect 2816 7588 2872 7590
rect 2896 7588 2952 7590
rect 2976 7588 3032 7590
rect 1916 7098 1972 7100
rect 1996 7098 2052 7100
rect 2076 7098 2132 7100
rect 2156 7098 2212 7100
rect 2236 7098 2292 7100
rect 1916 7046 1918 7098
rect 1918 7046 1970 7098
rect 1970 7046 1972 7098
rect 1996 7046 2034 7098
rect 2034 7046 2046 7098
rect 2046 7046 2052 7098
rect 2076 7046 2098 7098
rect 2098 7046 2110 7098
rect 2110 7046 2132 7098
rect 2156 7046 2162 7098
rect 2162 7046 2174 7098
rect 2174 7046 2212 7098
rect 2236 7046 2238 7098
rect 2238 7046 2290 7098
rect 2290 7046 2292 7098
rect 1916 7044 1972 7046
rect 1996 7044 2052 7046
rect 2076 7044 2132 7046
rect 2156 7044 2212 7046
rect 2236 7044 2292 7046
rect 1306 6568 1362 6624
rect 2656 6554 2712 6556
rect 2736 6554 2792 6556
rect 2816 6554 2872 6556
rect 2896 6554 2952 6556
rect 2976 6554 3032 6556
rect 2656 6502 2658 6554
rect 2658 6502 2710 6554
rect 2710 6502 2712 6554
rect 2736 6502 2774 6554
rect 2774 6502 2786 6554
rect 2786 6502 2792 6554
rect 2816 6502 2838 6554
rect 2838 6502 2850 6554
rect 2850 6502 2872 6554
rect 2896 6502 2902 6554
rect 2902 6502 2914 6554
rect 2914 6502 2952 6554
rect 2976 6502 2978 6554
rect 2978 6502 3030 6554
rect 3030 6502 3032 6554
rect 2656 6500 2712 6502
rect 2736 6500 2792 6502
rect 2816 6500 2872 6502
rect 2896 6500 2952 6502
rect 2976 6500 3032 6502
rect 1398 5516 1400 5536
rect 1400 5516 1452 5536
rect 1452 5516 1454 5536
rect 1398 5480 1454 5516
rect 846 4528 902 4584
rect 1916 6010 1972 6012
rect 1996 6010 2052 6012
rect 2076 6010 2132 6012
rect 2156 6010 2212 6012
rect 2236 6010 2292 6012
rect 1916 5958 1918 6010
rect 1918 5958 1970 6010
rect 1970 5958 1972 6010
rect 1996 5958 2034 6010
rect 2034 5958 2046 6010
rect 2046 5958 2052 6010
rect 2076 5958 2098 6010
rect 2098 5958 2110 6010
rect 2110 5958 2132 6010
rect 2156 5958 2162 6010
rect 2162 5958 2174 6010
rect 2174 5958 2212 6010
rect 2236 5958 2238 6010
rect 2238 5958 2290 6010
rect 2290 5958 2292 6010
rect 1916 5956 1972 5958
rect 1996 5956 2052 5958
rect 2076 5956 2132 5958
rect 2156 5956 2212 5958
rect 2236 5956 2292 5958
rect 1916 4922 1972 4924
rect 1996 4922 2052 4924
rect 2076 4922 2132 4924
rect 2156 4922 2212 4924
rect 2236 4922 2292 4924
rect 1916 4870 1918 4922
rect 1918 4870 1970 4922
rect 1970 4870 1972 4922
rect 1996 4870 2034 4922
rect 2034 4870 2046 4922
rect 2046 4870 2052 4922
rect 2076 4870 2098 4922
rect 2098 4870 2110 4922
rect 2110 4870 2132 4922
rect 2156 4870 2162 4922
rect 2162 4870 2174 4922
rect 2174 4870 2212 4922
rect 2236 4870 2238 4922
rect 2238 4870 2290 4922
rect 2290 4870 2292 4922
rect 1916 4868 1972 4870
rect 1996 4868 2052 4870
rect 2076 4868 2132 4870
rect 2156 4868 2212 4870
rect 2236 4868 2292 4870
rect 2656 5466 2712 5468
rect 2736 5466 2792 5468
rect 2816 5466 2872 5468
rect 2896 5466 2952 5468
rect 2976 5466 3032 5468
rect 2656 5414 2658 5466
rect 2658 5414 2710 5466
rect 2710 5414 2712 5466
rect 2736 5414 2774 5466
rect 2774 5414 2786 5466
rect 2786 5414 2792 5466
rect 2816 5414 2838 5466
rect 2838 5414 2850 5466
rect 2850 5414 2872 5466
rect 2896 5414 2902 5466
rect 2902 5414 2914 5466
rect 2914 5414 2952 5466
rect 2976 5414 2978 5466
rect 2978 5414 3030 5466
rect 3030 5414 3032 5466
rect 2656 5412 2712 5414
rect 2736 5412 2792 5414
rect 2816 5412 2872 5414
rect 2896 5412 2952 5414
rect 2976 5412 3032 5414
rect 846 3440 902 3496
rect 1916 3834 1972 3836
rect 1996 3834 2052 3836
rect 2076 3834 2132 3836
rect 2156 3834 2212 3836
rect 2236 3834 2292 3836
rect 1916 3782 1918 3834
rect 1918 3782 1970 3834
rect 1970 3782 1972 3834
rect 1996 3782 2034 3834
rect 2034 3782 2046 3834
rect 2046 3782 2052 3834
rect 2076 3782 2098 3834
rect 2098 3782 2110 3834
rect 2110 3782 2132 3834
rect 2156 3782 2162 3834
rect 2162 3782 2174 3834
rect 2174 3782 2212 3834
rect 2236 3782 2238 3834
rect 2238 3782 2290 3834
rect 2290 3782 2292 3834
rect 1916 3780 1972 3782
rect 1996 3780 2052 3782
rect 2076 3780 2132 3782
rect 2156 3780 2212 3782
rect 2236 3780 2292 3782
rect 2656 4378 2712 4380
rect 2736 4378 2792 4380
rect 2816 4378 2872 4380
rect 2896 4378 2952 4380
rect 2976 4378 3032 4380
rect 2656 4326 2658 4378
rect 2658 4326 2710 4378
rect 2710 4326 2712 4378
rect 2736 4326 2774 4378
rect 2774 4326 2786 4378
rect 2786 4326 2792 4378
rect 2816 4326 2838 4378
rect 2838 4326 2850 4378
rect 2850 4326 2872 4378
rect 2896 4326 2902 4378
rect 2902 4326 2914 4378
rect 2914 4326 2952 4378
rect 2976 4326 2978 4378
rect 2978 4326 3030 4378
rect 3030 4326 3032 4378
rect 2656 4324 2712 4326
rect 2736 4324 2792 4326
rect 2816 4324 2872 4326
rect 2896 4324 2952 4326
rect 2976 4324 3032 4326
rect 2656 3290 2712 3292
rect 2736 3290 2792 3292
rect 2816 3290 2872 3292
rect 2896 3290 2952 3292
rect 2976 3290 3032 3292
rect 2656 3238 2658 3290
rect 2658 3238 2710 3290
rect 2710 3238 2712 3290
rect 2736 3238 2774 3290
rect 2774 3238 2786 3290
rect 2786 3238 2792 3290
rect 2816 3238 2838 3290
rect 2838 3238 2850 3290
rect 2850 3238 2872 3290
rect 2896 3238 2902 3290
rect 2902 3238 2914 3290
rect 2914 3238 2952 3290
rect 2976 3238 2978 3290
rect 2978 3238 3030 3290
rect 3030 3238 3032 3290
rect 2656 3236 2712 3238
rect 2736 3236 2792 3238
rect 2816 3236 2872 3238
rect 2896 3236 2952 3238
rect 2976 3236 3032 3238
rect 8656 18522 8712 18524
rect 8736 18522 8792 18524
rect 8816 18522 8872 18524
rect 8896 18522 8952 18524
rect 8976 18522 9032 18524
rect 8656 18470 8658 18522
rect 8658 18470 8710 18522
rect 8710 18470 8712 18522
rect 8736 18470 8774 18522
rect 8774 18470 8786 18522
rect 8786 18470 8792 18522
rect 8816 18470 8838 18522
rect 8838 18470 8850 18522
rect 8850 18470 8872 18522
rect 8896 18470 8902 18522
rect 8902 18470 8914 18522
rect 8914 18470 8952 18522
rect 8976 18470 8978 18522
rect 8978 18470 9030 18522
rect 9030 18470 9032 18522
rect 8656 18468 8712 18470
rect 8736 18468 8792 18470
rect 8816 18468 8872 18470
rect 8896 18468 8952 18470
rect 8976 18468 9032 18470
rect 14656 18522 14712 18524
rect 14736 18522 14792 18524
rect 14816 18522 14872 18524
rect 14896 18522 14952 18524
rect 14976 18522 15032 18524
rect 14656 18470 14658 18522
rect 14658 18470 14710 18522
rect 14710 18470 14712 18522
rect 14736 18470 14774 18522
rect 14774 18470 14786 18522
rect 14786 18470 14792 18522
rect 14816 18470 14838 18522
rect 14838 18470 14850 18522
rect 14850 18470 14872 18522
rect 14896 18470 14902 18522
rect 14902 18470 14914 18522
rect 14914 18470 14952 18522
rect 14976 18470 14978 18522
rect 14978 18470 15030 18522
rect 15030 18470 15032 18522
rect 14656 18468 14712 18470
rect 14736 18468 14792 18470
rect 14816 18468 14872 18470
rect 14896 18468 14952 18470
rect 14976 18468 15032 18470
rect 7916 17978 7972 17980
rect 7996 17978 8052 17980
rect 8076 17978 8132 17980
rect 8156 17978 8212 17980
rect 8236 17978 8292 17980
rect 7916 17926 7918 17978
rect 7918 17926 7970 17978
rect 7970 17926 7972 17978
rect 7996 17926 8034 17978
rect 8034 17926 8046 17978
rect 8046 17926 8052 17978
rect 8076 17926 8098 17978
rect 8098 17926 8110 17978
rect 8110 17926 8132 17978
rect 8156 17926 8162 17978
rect 8162 17926 8174 17978
rect 8174 17926 8212 17978
rect 8236 17926 8238 17978
rect 8238 17926 8290 17978
rect 8290 17926 8292 17978
rect 7916 17924 7972 17926
rect 7996 17924 8052 17926
rect 8076 17924 8132 17926
rect 8156 17924 8212 17926
rect 8236 17924 8292 17926
rect 8656 17434 8712 17436
rect 8736 17434 8792 17436
rect 8816 17434 8872 17436
rect 8896 17434 8952 17436
rect 8976 17434 9032 17436
rect 8656 17382 8658 17434
rect 8658 17382 8710 17434
rect 8710 17382 8712 17434
rect 8736 17382 8774 17434
rect 8774 17382 8786 17434
rect 8786 17382 8792 17434
rect 8816 17382 8838 17434
rect 8838 17382 8850 17434
rect 8850 17382 8872 17434
rect 8896 17382 8902 17434
rect 8902 17382 8914 17434
rect 8914 17382 8952 17434
rect 8976 17382 8978 17434
rect 8978 17382 9030 17434
rect 9030 17382 9032 17434
rect 8656 17380 8712 17382
rect 8736 17380 8792 17382
rect 8816 17380 8872 17382
rect 8896 17380 8952 17382
rect 8976 17380 9032 17382
rect 7916 16890 7972 16892
rect 7996 16890 8052 16892
rect 8076 16890 8132 16892
rect 8156 16890 8212 16892
rect 8236 16890 8292 16892
rect 7916 16838 7918 16890
rect 7918 16838 7970 16890
rect 7970 16838 7972 16890
rect 7996 16838 8034 16890
rect 8034 16838 8046 16890
rect 8046 16838 8052 16890
rect 8076 16838 8098 16890
rect 8098 16838 8110 16890
rect 8110 16838 8132 16890
rect 8156 16838 8162 16890
rect 8162 16838 8174 16890
rect 8174 16838 8212 16890
rect 8236 16838 8238 16890
rect 8238 16838 8290 16890
rect 8290 16838 8292 16890
rect 7916 16836 7972 16838
rect 7996 16836 8052 16838
rect 8076 16836 8132 16838
rect 8156 16836 8212 16838
rect 8236 16836 8292 16838
rect 8656 16346 8712 16348
rect 8736 16346 8792 16348
rect 8816 16346 8872 16348
rect 8896 16346 8952 16348
rect 8976 16346 9032 16348
rect 8656 16294 8658 16346
rect 8658 16294 8710 16346
rect 8710 16294 8712 16346
rect 8736 16294 8774 16346
rect 8774 16294 8786 16346
rect 8786 16294 8792 16346
rect 8816 16294 8838 16346
rect 8838 16294 8850 16346
rect 8850 16294 8872 16346
rect 8896 16294 8902 16346
rect 8902 16294 8914 16346
rect 8914 16294 8952 16346
rect 8976 16294 8978 16346
rect 8978 16294 9030 16346
rect 9030 16294 9032 16346
rect 8656 16292 8712 16294
rect 8736 16292 8792 16294
rect 8816 16292 8872 16294
rect 8896 16292 8952 16294
rect 8976 16292 9032 16294
rect 7916 15802 7972 15804
rect 7996 15802 8052 15804
rect 8076 15802 8132 15804
rect 8156 15802 8212 15804
rect 8236 15802 8292 15804
rect 7916 15750 7918 15802
rect 7918 15750 7970 15802
rect 7970 15750 7972 15802
rect 7996 15750 8034 15802
rect 8034 15750 8046 15802
rect 8046 15750 8052 15802
rect 8076 15750 8098 15802
rect 8098 15750 8110 15802
rect 8110 15750 8132 15802
rect 8156 15750 8162 15802
rect 8162 15750 8174 15802
rect 8174 15750 8212 15802
rect 8236 15750 8238 15802
rect 8238 15750 8290 15802
rect 8290 15750 8292 15802
rect 7916 15748 7972 15750
rect 7996 15748 8052 15750
rect 8076 15748 8132 15750
rect 8156 15748 8212 15750
rect 8236 15748 8292 15750
rect 8656 15258 8712 15260
rect 8736 15258 8792 15260
rect 8816 15258 8872 15260
rect 8896 15258 8952 15260
rect 8976 15258 9032 15260
rect 8656 15206 8658 15258
rect 8658 15206 8710 15258
rect 8710 15206 8712 15258
rect 8736 15206 8774 15258
rect 8774 15206 8786 15258
rect 8786 15206 8792 15258
rect 8816 15206 8838 15258
rect 8838 15206 8850 15258
rect 8850 15206 8872 15258
rect 8896 15206 8902 15258
rect 8902 15206 8914 15258
rect 8914 15206 8952 15258
rect 8976 15206 8978 15258
rect 8978 15206 9030 15258
rect 9030 15206 9032 15258
rect 8656 15204 8712 15206
rect 8736 15204 8792 15206
rect 8816 15204 8872 15206
rect 8896 15204 8952 15206
rect 8976 15204 9032 15206
rect 7916 14714 7972 14716
rect 7996 14714 8052 14716
rect 8076 14714 8132 14716
rect 8156 14714 8212 14716
rect 8236 14714 8292 14716
rect 7916 14662 7918 14714
rect 7918 14662 7970 14714
rect 7970 14662 7972 14714
rect 7996 14662 8034 14714
rect 8034 14662 8046 14714
rect 8046 14662 8052 14714
rect 8076 14662 8098 14714
rect 8098 14662 8110 14714
rect 8110 14662 8132 14714
rect 8156 14662 8162 14714
rect 8162 14662 8174 14714
rect 8174 14662 8212 14714
rect 8236 14662 8238 14714
rect 8238 14662 8290 14714
rect 8290 14662 8292 14714
rect 7916 14660 7972 14662
rect 7996 14660 8052 14662
rect 8076 14660 8132 14662
rect 8156 14660 8212 14662
rect 8236 14660 8292 14662
rect 8656 14170 8712 14172
rect 8736 14170 8792 14172
rect 8816 14170 8872 14172
rect 8896 14170 8952 14172
rect 8976 14170 9032 14172
rect 8656 14118 8658 14170
rect 8658 14118 8710 14170
rect 8710 14118 8712 14170
rect 8736 14118 8774 14170
rect 8774 14118 8786 14170
rect 8786 14118 8792 14170
rect 8816 14118 8838 14170
rect 8838 14118 8850 14170
rect 8850 14118 8872 14170
rect 8896 14118 8902 14170
rect 8902 14118 8914 14170
rect 8914 14118 8952 14170
rect 8976 14118 8978 14170
rect 8978 14118 9030 14170
rect 9030 14118 9032 14170
rect 8656 14116 8712 14118
rect 8736 14116 8792 14118
rect 8816 14116 8872 14118
rect 8896 14116 8952 14118
rect 8976 14116 9032 14118
rect 7916 13626 7972 13628
rect 7996 13626 8052 13628
rect 8076 13626 8132 13628
rect 8156 13626 8212 13628
rect 8236 13626 8292 13628
rect 7916 13574 7918 13626
rect 7918 13574 7970 13626
rect 7970 13574 7972 13626
rect 7996 13574 8034 13626
rect 8034 13574 8046 13626
rect 8046 13574 8052 13626
rect 8076 13574 8098 13626
rect 8098 13574 8110 13626
rect 8110 13574 8132 13626
rect 8156 13574 8162 13626
rect 8162 13574 8174 13626
rect 8174 13574 8212 13626
rect 8236 13574 8238 13626
rect 8238 13574 8290 13626
rect 8290 13574 8292 13626
rect 7916 13572 7972 13574
rect 7996 13572 8052 13574
rect 8076 13572 8132 13574
rect 8156 13572 8212 13574
rect 8236 13572 8292 13574
rect 8656 13082 8712 13084
rect 8736 13082 8792 13084
rect 8816 13082 8872 13084
rect 8896 13082 8952 13084
rect 8976 13082 9032 13084
rect 8656 13030 8658 13082
rect 8658 13030 8710 13082
rect 8710 13030 8712 13082
rect 8736 13030 8774 13082
rect 8774 13030 8786 13082
rect 8786 13030 8792 13082
rect 8816 13030 8838 13082
rect 8838 13030 8850 13082
rect 8850 13030 8872 13082
rect 8896 13030 8902 13082
rect 8902 13030 8914 13082
rect 8914 13030 8952 13082
rect 8976 13030 8978 13082
rect 8978 13030 9030 13082
rect 9030 13030 9032 13082
rect 8656 13028 8712 13030
rect 8736 13028 8792 13030
rect 8816 13028 8872 13030
rect 8896 13028 8952 13030
rect 8976 13028 9032 13030
rect 7916 12538 7972 12540
rect 7996 12538 8052 12540
rect 8076 12538 8132 12540
rect 8156 12538 8212 12540
rect 8236 12538 8292 12540
rect 7916 12486 7918 12538
rect 7918 12486 7970 12538
rect 7970 12486 7972 12538
rect 7996 12486 8034 12538
rect 8034 12486 8046 12538
rect 8046 12486 8052 12538
rect 8076 12486 8098 12538
rect 8098 12486 8110 12538
rect 8110 12486 8132 12538
rect 8156 12486 8162 12538
rect 8162 12486 8174 12538
rect 8174 12486 8212 12538
rect 8236 12486 8238 12538
rect 8238 12486 8290 12538
rect 8290 12486 8292 12538
rect 7916 12484 7972 12486
rect 7996 12484 8052 12486
rect 8076 12484 8132 12486
rect 8156 12484 8212 12486
rect 8236 12484 8292 12486
rect 8656 11994 8712 11996
rect 8736 11994 8792 11996
rect 8816 11994 8872 11996
rect 8896 11994 8952 11996
rect 8976 11994 9032 11996
rect 8656 11942 8658 11994
rect 8658 11942 8710 11994
rect 8710 11942 8712 11994
rect 8736 11942 8774 11994
rect 8774 11942 8786 11994
rect 8786 11942 8792 11994
rect 8816 11942 8838 11994
rect 8838 11942 8850 11994
rect 8850 11942 8872 11994
rect 8896 11942 8902 11994
rect 8902 11942 8914 11994
rect 8914 11942 8952 11994
rect 8976 11942 8978 11994
rect 8978 11942 9030 11994
rect 9030 11942 9032 11994
rect 8656 11940 8712 11942
rect 8736 11940 8792 11942
rect 8816 11940 8872 11942
rect 8896 11940 8952 11942
rect 8976 11940 9032 11942
rect 7916 11450 7972 11452
rect 7996 11450 8052 11452
rect 8076 11450 8132 11452
rect 8156 11450 8212 11452
rect 8236 11450 8292 11452
rect 7916 11398 7918 11450
rect 7918 11398 7970 11450
rect 7970 11398 7972 11450
rect 7996 11398 8034 11450
rect 8034 11398 8046 11450
rect 8046 11398 8052 11450
rect 8076 11398 8098 11450
rect 8098 11398 8110 11450
rect 8110 11398 8132 11450
rect 8156 11398 8162 11450
rect 8162 11398 8174 11450
rect 8174 11398 8212 11450
rect 8236 11398 8238 11450
rect 8238 11398 8290 11450
rect 8290 11398 8292 11450
rect 7916 11396 7972 11398
rect 7996 11396 8052 11398
rect 8076 11396 8132 11398
rect 8156 11396 8212 11398
rect 8236 11396 8292 11398
rect 6734 6316 6790 6352
rect 6734 6296 6736 6316
rect 6736 6296 6788 6316
rect 6788 6296 6790 6316
rect 7916 10362 7972 10364
rect 7996 10362 8052 10364
rect 8076 10362 8132 10364
rect 8156 10362 8212 10364
rect 8236 10362 8292 10364
rect 7916 10310 7918 10362
rect 7918 10310 7970 10362
rect 7970 10310 7972 10362
rect 7996 10310 8034 10362
rect 8034 10310 8046 10362
rect 8046 10310 8052 10362
rect 8076 10310 8098 10362
rect 8098 10310 8110 10362
rect 8110 10310 8132 10362
rect 8156 10310 8162 10362
rect 8162 10310 8174 10362
rect 8174 10310 8212 10362
rect 8236 10310 8238 10362
rect 8238 10310 8290 10362
rect 8290 10310 8292 10362
rect 7916 10308 7972 10310
rect 7996 10308 8052 10310
rect 8076 10308 8132 10310
rect 8156 10308 8212 10310
rect 8236 10308 8292 10310
rect 7916 9274 7972 9276
rect 7996 9274 8052 9276
rect 8076 9274 8132 9276
rect 8156 9274 8212 9276
rect 8236 9274 8292 9276
rect 7916 9222 7918 9274
rect 7918 9222 7970 9274
rect 7970 9222 7972 9274
rect 7996 9222 8034 9274
rect 8034 9222 8046 9274
rect 8046 9222 8052 9274
rect 8076 9222 8098 9274
rect 8098 9222 8110 9274
rect 8110 9222 8132 9274
rect 8156 9222 8162 9274
rect 8162 9222 8174 9274
rect 8174 9222 8212 9274
rect 8236 9222 8238 9274
rect 8238 9222 8290 9274
rect 8290 9222 8292 9274
rect 7916 9220 7972 9222
rect 7996 9220 8052 9222
rect 8076 9220 8132 9222
rect 8156 9220 8212 9222
rect 8236 9220 8292 9222
rect 8656 10906 8712 10908
rect 8736 10906 8792 10908
rect 8816 10906 8872 10908
rect 8896 10906 8952 10908
rect 8976 10906 9032 10908
rect 8656 10854 8658 10906
rect 8658 10854 8710 10906
rect 8710 10854 8712 10906
rect 8736 10854 8774 10906
rect 8774 10854 8786 10906
rect 8786 10854 8792 10906
rect 8816 10854 8838 10906
rect 8838 10854 8850 10906
rect 8850 10854 8872 10906
rect 8896 10854 8902 10906
rect 8902 10854 8914 10906
rect 8914 10854 8952 10906
rect 8976 10854 8978 10906
rect 8978 10854 9030 10906
rect 9030 10854 9032 10906
rect 8656 10852 8712 10854
rect 8736 10852 8792 10854
rect 8816 10852 8872 10854
rect 8896 10852 8952 10854
rect 8976 10852 9032 10854
rect 8656 9818 8712 9820
rect 8736 9818 8792 9820
rect 8816 9818 8872 9820
rect 8896 9818 8952 9820
rect 8976 9818 9032 9820
rect 8656 9766 8658 9818
rect 8658 9766 8710 9818
rect 8710 9766 8712 9818
rect 8736 9766 8774 9818
rect 8774 9766 8786 9818
rect 8786 9766 8792 9818
rect 8816 9766 8838 9818
rect 8838 9766 8850 9818
rect 8850 9766 8872 9818
rect 8896 9766 8902 9818
rect 8902 9766 8914 9818
rect 8914 9766 8952 9818
rect 8976 9766 8978 9818
rect 8978 9766 9030 9818
rect 9030 9766 9032 9818
rect 8656 9764 8712 9766
rect 8736 9764 8792 9766
rect 8816 9764 8872 9766
rect 8896 9764 8952 9766
rect 8976 9764 9032 9766
rect 8656 8730 8712 8732
rect 8736 8730 8792 8732
rect 8816 8730 8872 8732
rect 8896 8730 8952 8732
rect 8976 8730 9032 8732
rect 8656 8678 8658 8730
rect 8658 8678 8710 8730
rect 8710 8678 8712 8730
rect 8736 8678 8774 8730
rect 8774 8678 8786 8730
rect 8786 8678 8792 8730
rect 8816 8678 8838 8730
rect 8838 8678 8850 8730
rect 8850 8678 8872 8730
rect 8896 8678 8902 8730
rect 8902 8678 8914 8730
rect 8914 8678 8952 8730
rect 8976 8678 8978 8730
rect 8978 8678 9030 8730
rect 9030 8678 9032 8730
rect 8656 8676 8712 8678
rect 8736 8676 8792 8678
rect 8816 8676 8872 8678
rect 8896 8676 8952 8678
rect 8976 8676 9032 8678
rect 7916 8186 7972 8188
rect 7996 8186 8052 8188
rect 8076 8186 8132 8188
rect 8156 8186 8212 8188
rect 8236 8186 8292 8188
rect 7916 8134 7918 8186
rect 7918 8134 7970 8186
rect 7970 8134 7972 8186
rect 7996 8134 8034 8186
rect 8034 8134 8046 8186
rect 8046 8134 8052 8186
rect 8076 8134 8098 8186
rect 8098 8134 8110 8186
rect 8110 8134 8132 8186
rect 8156 8134 8162 8186
rect 8162 8134 8174 8186
rect 8174 8134 8212 8186
rect 8236 8134 8238 8186
rect 8238 8134 8290 8186
rect 8290 8134 8292 8186
rect 7916 8132 7972 8134
rect 7996 8132 8052 8134
rect 8076 8132 8132 8134
rect 8156 8132 8212 8134
rect 8236 8132 8292 8134
rect 8656 7642 8712 7644
rect 8736 7642 8792 7644
rect 8816 7642 8872 7644
rect 8896 7642 8952 7644
rect 8976 7642 9032 7644
rect 8656 7590 8658 7642
rect 8658 7590 8710 7642
rect 8710 7590 8712 7642
rect 8736 7590 8774 7642
rect 8774 7590 8786 7642
rect 8786 7590 8792 7642
rect 8816 7590 8838 7642
rect 8838 7590 8850 7642
rect 8850 7590 8872 7642
rect 8896 7590 8902 7642
rect 8902 7590 8914 7642
rect 8914 7590 8952 7642
rect 8976 7590 8978 7642
rect 8978 7590 9030 7642
rect 9030 7590 9032 7642
rect 8656 7588 8712 7590
rect 8736 7588 8792 7590
rect 8816 7588 8872 7590
rect 8896 7588 8952 7590
rect 8976 7588 9032 7590
rect 7916 7098 7972 7100
rect 7996 7098 8052 7100
rect 8076 7098 8132 7100
rect 8156 7098 8212 7100
rect 8236 7098 8292 7100
rect 7916 7046 7918 7098
rect 7918 7046 7970 7098
rect 7970 7046 7972 7098
rect 7996 7046 8034 7098
rect 8034 7046 8046 7098
rect 8046 7046 8052 7098
rect 8076 7046 8098 7098
rect 8098 7046 8110 7098
rect 8110 7046 8132 7098
rect 8156 7046 8162 7098
rect 8162 7046 8174 7098
rect 8174 7046 8212 7098
rect 8236 7046 8238 7098
rect 8238 7046 8290 7098
rect 8290 7046 8292 7098
rect 7916 7044 7972 7046
rect 7996 7044 8052 7046
rect 8076 7044 8132 7046
rect 8156 7044 8212 7046
rect 8236 7044 8292 7046
rect 7838 6840 7894 6896
rect 1916 2746 1972 2748
rect 1996 2746 2052 2748
rect 2076 2746 2132 2748
rect 2156 2746 2212 2748
rect 2236 2746 2292 2748
rect 1916 2694 1918 2746
rect 1918 2694 1970 2746
rect 1970 2694 1972 2746
rect 1996 2694 2034 2746
rect 2034 2694 2046 2746
rect 2046 2694 2052 2746
rect 2076 2694 2098 2746
rect 2098 2694 2110 2746
rect 2110 2694 2132 2746
rect 2156 2694 2162 2746
rect 2162 2694 2174 2746
rect 2174 2694 2212 2746
rect 2236 2694 2238 2746
rect 2238 2694 2290 2746
rect 2290 2694 2292 2746
rect 1916 2692 1972 2694
rect 1996 2692 2052 2694
rect 2076 2692 2132 2694
rect 2156 2692 2212 2694
rect 2236 2692 2292 2694
rect 7562 6724 7618 6760
rect 7562 6704 7564 6724
rect 7564 6704 7616 6724
rect 7616 6704 7618 6724
rect 9402 6740 9404 6760
rect 9404 6740 9456 6760
rect 9456 6740 9458 6760
rect 7916 6010 7972 6012
rect 7996 6010 8052 6012
rect 8076 6010 8132 6012
rect 8156 6010 8212 6012
rect 8236 6010 8292 6012
rect 7916 5958 7918 6010
rect 7918 5958 7970 6010
rect 7970 5958 7972 6010
rect 7996 5958 8034 6010
rect 8034 5958 8046 6010
rect 8046 5958 8052 6010
rect 8076 5958 8098 6010
rect 8098 5958 8110 6010
rect 8110 5958 8132 6010
rect 8156 5958 8162 6010
rect 8162 5958 8174 6010
rect 8174 5958 8212 6010
rect 8236 5958 8238 6010
rect 8238 5958 8290 6010
rect 8290 5958 8292 6010
rect 7916 5956 7972 5958
rect 7996 5956 8052 5958
rect 8076 5956 8132 5958
rect 8156 5956 8212 5958
rect 8236 5956 8292 5958
rect 8656 6554 8712 6556
rect 8736 6554 8792 6556
rect 8816 6554 8872 6556
rect 8896 6554 8952 6556
rect 8976 6554 9032 6556
rect 8656 6502 8658 6554
rect 8658 6502 8710 6554
rect 8710 6502 8712 6554
rect 8736 6502 8774 6554
rect 8774 6502 8786 6554
rect 8786 6502 8792 6554
rect 8816 6502 8838 6554
rect 8838 6502 8850 6554
rect 8850 6502 8872 6554
rect 8896 6502 8902 6554
rect 8902 6502 8914 6554
rect 8914 6502 8952 6554
rect 8976 6502 8978 6554
rect 8978 6502 9030 6554
rect 9030 6502 9032 6554
rect 8656 6500 8712 6502
rect 8736 6500 8792 6502
rect 8816 6500 8872 6502
rect 8896 6500 8952 6502
rect 8976 6500 9032 6502
rect 9402 6704 9458 6740
rect 7916 4922 7972 4924
rect 7996 4922 8052 4924
rect 8076 4922 8132 4924
rect 8156 4922 8212 4924
rect 8236 4922 8292 4924
rect 7916 4870 7918 4922
rect 7918 4870 7970 4922
rect 7970 4870 7972 4922
rect 7996 4870 8034 4922
rect 8034 4870 8046 4922
rect 8046 4870 8052 4922
rect 8076 4870 8098 4922
rect 8098 4870 8110 4922
rect 8110 4870 8132 4922
rect 8156 4870 8162 4922
rect 8162 4870 8174 4922
rect 8174 4870 8212 4922
rect 8236 4870 8238 4922
rect 8238 4870 8290 4922
rect 8290 4870 8292 4922
rect 7916 4868 7972 4870
rect 7996 4868 8052 4870
rect 8076 4868 8132 4870
rect 8156 4868 8212 4870
rect 8236 4868 8292 4870
rect 7916 3834 7972 3836
rect 7996 3834 8052 3836
rect 8076 3834 8132 3836
rect 8156 3834 8212 3836
rect 8236 3834 8292 3836
rect 7916 3782 7918 3834
rect 7918 3782 7970 3834
rect 7970 3782 7972 3834
rect 7996 3782 8034 3834
rect 8034 3782 8046 3834
rect 8046 3782 8052 3834
rect 8076 3782 8098 3834
rect 8098 3782 8110 3834
rect 8110 3782 8132 3834
rect 8156 3782 8162 3834
rect 8162 3782 8174 3834
rect 8174 3782 8212 3834
rect 8236 3782 8238 3834
rect 8238 3782 8290 3834
rect 8290 3782 8292 3834
rect 7916 3780 7972 3782
rect 7996 3780 8052 3782
rect 8076 3780 8132 3782
rect 8156 3780 8212 3782
rect 8236 3780 8292 3782
rect 8656 5466 8712 5468
rect 8736 5466 8792 5468
rect 8816 5466 8872 5468
rect 8896 5466 8952 5468
rect 8976 5466 9032 5468
rect 8656 5414 8658 5466
rect 8658 5414 8710 5466
rect 8710 5414 8712 5466
rect 8736 5414 8774 5466
rect 8774 5414 8786 5466
rect 8786 5414 8792 5466
rect 8816 5414 8838 5466
rect 8838 5414 8850 5466
rect 8850 5414 8872 5466
rect 8896 5414 8902 5466
rect 8902 5414 8914 5466
rect 8914 5414 8952 5466
rect 8976 5414 8978 5466
rect 8978 5414 9030 5466
rect 9030 5414 9032 5466
rect 8656 5412 8712 5414
rect 8736 5412 8792 5414
rect 8816 5412 8872 5414
rect 8896 5412 8952 5414
rect 8976 5412 9032 5414
rect 10690 6160 10746 6216
rect 8656 4378 8712 4380
rect 8736 4378 8792 4380
rect 8816 4378 8872 4380
rect 8896 4378 8952 4380
rect 8976 4378 9032 4380
rect 8656 4326 8658 4378
rect 8658 4326 8710 4378
rect 8710 4326 8712 4378
rect 8736 4326 8774 4378
rect 8774 4326 8786 4378
rect 8786 4326 8792 4378
rect 8816 4326 8838 4378
rect 8838 4326 8850 4378
rect 8850 4326 8872 4378
rect 8896 4326 8902 4378
rect 8902 4326 8914 4378
rect 8914 4326 8952 4378
rect 8976 4326 8978 4378
rect 8978 4326 9030 4378
rect 9030 4326 9032 4378
rect 8656 4324 8712 4326
rect 8736 4324 8792 4326
rect 8816 4324 8872 4326
rect 8896 4324 8952 4326
rect 8976 4324 9032 4326
rect 9770 3984 9826 4040
rect 8656 3290 8712 3292
rect 8736 3290 8792 3292
rect 8816 3290 8872 3292
rect 8896 3290 8952 3292
rect 8976 3290 9032 3292
rect 8656 3238 8658 3290
rect 8658 3238 8710 3290
rect 8710 3238 8712 3290
rect 8736 3238 8774 3290
rect 8774 3238 8786 3290
rect 8786 3238 8792 3290
rect 8816 3238 8838 3290
rect 8838 3238 8850 3290
rect 8850 3238 8872 3290
rect 8896 3238 8902 3290
rect 8902 3238 8914 3290
rect 8914 3238 8952 3290
rect 8976 3238 8978 3290
rect 8978 3238 9030 3290
rect 9030 3238 9032 3290
rect 8656 3236 8712 3238
rect 8736 3236 8792 3238
rect 8816 3236 8872 3238
rect 8896 3236 8952 3238
rect 8976 3236 9032 3238
rect 7916 2746 7972 2748
rect 7996 2746 8052 2748
rect 8076 2746 8132 2748
rect 8156 2746 8212 2748
rect 8236 2746 8292 2748
rect 7916 2694 7918 2746
rect 7918 2694 7970 2746
rect 7970 2694 7972 2746
rect 7996 2694 8034 2746
rect 8034 2694 8046 2746
rect 8046 2694 8052 2746
rect 8076 2694 8098 2746
rect 8098 2694 8110 2746
rect 8110 2694 8132 2746
rect 8156 2694 8162 2746
rect 8162 2694 8174 2746
rect 8174 2694 8212 2746
rect 8236 2694 8238 2746
rect 8238 2694 8290 2746
rect 8290 2694 8292 2746
rect 7916 2692 7972 2694
rect 7996 2692 8052 2694
rect 8076 2692 8132 2694
rect 8156 2692 8212 2694
rect 8236 2692 8292 2694
rect 12438 18028 12440 18048
rect 12440 18028 12492 18048
rect 12492 18028 12494 18048
rect 12438 17992 12494 18028
rect 13916 17978 13972 17980
rect 13996 17978 14052 17980
rect 14076 17978 14132 17980
rect 14156 17978 14212 17980
rect 14236 17978 14292 17980
rect 13916 17926 13918 17978
rect 13918 17926 13970 17978
rect 13970 17926 13972 17978
rect 13996 17926 14034 17978
rect 14034 17926 14046 17978
rect 14046 17926 14052 17978
rect 14076 17926 14098 17978
rect 14098 17926 14110 17978
rect 14110 17926 14132 17978
rect 14156 17926 14162 17978
rect 14162 17926 14174 17978
rect 14174 17926 14212 17978
rect 14236 17926 14238 17978
rect 14238 17926 14290 17978
rect 14290 17926 14292 17978
rect 13916 17924 13972 17926
rect 13996 17924 14052 17926
rect 14076 17924 14132 17926
rect 14156 17924 14212 17926
rect 14236 17924 14292 17926
rect 12070 15544 12126 15600
rect 14656 17434 14712 17436
rect 14736 17434 14792 17436
rect 14816 17434 14872 17436
rect 14896 17434 14952 17436
rect 14976 17434 15032 17436
rect 14656 17382 14658 17434
rect 14658 17382 14710 17434
rect 14710 17382 14712 17434
rect 14736 17382 14774 17434
rect 14774 17382 14786 17434
rect 14786 17382 14792 17434
rect 14816 17382 14838 17434
rect 14838 17382 14850 17434
rect 14850 17382 14872 17434
rect 14896 17382 14902 17434
rect 14902 17382 14914 17434
rect 14914 17382 14952 17434
rect 14976 17382 14978 17434
rect 14978 17382 15030 17434
rect 15030 17382 15032 17434
rect 14656 17380 14712 17382
rect 14736 17380 14792 17382
rect 14816 17380 14872 17382
rect 14896 17380 14952 17382
rect 14976 17380 15032 17382
rect 13916 16890 13972 16892
rect 13996 16890 14052 16892
rect 14076 16890 14132 16892
rect 14156 16890 14212 16892
rect 14236 16890 14292 16892
rect 13916 16838 13918 16890
rect 13918 16838 13970 16890
rect 13970 16838 13972 16890
rect 13996 16838 14034 16890
rect 14034 16838 14046 16890
rect 14046 16838 14052 16890
rect 14076 16838 14098 16890
rect 14098 16838 14110 16890
rect 14110 16838 14132 16890
rect 14156 16838 14162 16890
rect 14162 16838 14174 16890
rect 14174 16838 14212 16890
rect 14236 16838 14238 16890
rect 14238 16838 14290 16890
rect 14290 16838 14292 16890
rect 13916 16836 13972 16838
rect 13996 16836 14052 16838
rect 14076 16836 14132 16838
rect 14156 16836 14212 16838
rect 14236 16836 14292 16838
rect 12714 15544 12770 15600
rect 14656 16346 14712 16348
rect 14736 16346 14792 16348
rect 14816 16346 14872 16348
rect 14896 16346 14952 16348
rect 14976 16346 15032 16348
rect 14656 16294 14658 16346
rect 14658 16294 14710 16346
rect 14710 16294 14712 16346
rect 14736 16294 14774 16346
rect 14774 16294 14786 16346
rect 14786 16294 14792 16346
rect 14816 16294 14838 16346
rect 14838 16294 14850 16346
rect 14850 16294 14872 16346
rect 14896 16294 14902 16346
rect 14902 16294 14914 16346
rect 14914 16294 14952 16346
rect 14976 16294 14978 16346
rect 14978 16294 15030 16346
rect 15030 16294 15032 16346
rect 14656 16292 14712 16294
rect 14736 16292 14792 16294
rect 14816 16292 14872 16294
rect 14896 16292 14952 16294
rect 14976 16292 15032 16294
rect 13916 15802 13972 15804
rect 13996 15802 14052 15804
rect 14076 15802 14132 15804
rect 14156 15802 14212 15804
rect 14236 15802 14292 15804
rect 13916 15750 13918 15802
rect 13918 15750 13970 15802
rect 13970 15750 13972 15802
rect 13996 15750 14034 15802
rect 14034 15750 14046 15802
rect 14046 15750 14052 15802
rect 14076 15750 14098 15802
rect 14098 15750 14110 15802
rect 14110 15750 14132 15802
rect 14156 15750 14162 15802
rect 14162 15750 14174 15802
rect 14174 15750 14212 15802
rect 14236 15750 14238 15802
rect 14238 15750 14290 15802
rect 14290 15750 14292 15802
rect 13916 15748 13972 15750
rect 13996 15748 14052 15750
rect 14076 15748 14132 15750
rect 14156 15748 14212 15750
rect 14236 15748 14292 15750
rect 13916 14714 13972 14716
rect 13996 14714 14052 14716
rect 14076 14714 14132 14716
rect 14156 14714 14212 14716
rect 14236 14714 14292 14716
rect 13916 14662 13918 14714
rect 13918 14662 13970 14714
rect 13970 14662 13972 14714
rect 13996 14662 14034 14714
rect 14034 14662 14046 14714
rect 14046 14662 14052 14714
rect 14076 14662 14098 14714
rect 14098 14662 14110 14714
rect 14110 14662 14132 14714
rect 14156 14662 14162 14714
rect 14162 14662 14174 14714
rect 14174 14662 14212 14714
rect 14236 14662 14238 14714
rect 14238 14662 14290 14714
rect 14290 14662 14292 14714
rect 13916 14660 13972 14662
rect 13996 14660 14052 14662
rect 14076 14660 14132 14662
rect 14156 14660 14212 14662
rect 14236 14660 14292 14662
rect 14656 15258 14712 15260
rect 14736 15258 14792 15260
rect 14816 15258 14872 15260
rect 14896 15258 14952 15260
rect 14976 15258 15032 15260
rect 14656 15206 14658 15258
rect 14658 15206 14710 15258
rect 14710 15206 14712 15258
rect 14736 15206 14774 15258
rect 14774 15206 14786 15258
rect 14786 15206 14792 15258
rect 14816 15206 14838 15258
rect 14838 15206 14850 15258
rect 14850 15206 14872 15258
rect 14896 15206 14902 15258
rect 14902 15206 14914 15258
rect 14914 15206 14952 15258
rect 14976 15206 14978 15258
rect 14978 15206 15030 15258
rect 15030 15206 15032 15258
rect 14656 15204 14712 15206
rect 14736 15204 14792 15206
rect 14816 15204 14872 15206
rect 14896 15204 14952 15206
rect 14976 15204 15032 15206
rect 14656 14170 14712 14172
rect 14736 14170 14792 14172
rect 14816 14170 14872 14172
rect 14896 14170 14952 14172
rect 14976 14170 15032 14172
rect 14656 14118 14658 14170
rect 14658 14118 14710 14170
rect 14710 14118 14712 14170
rect 14736 14118 14774 14170
rect 14774 14118 14786 14170
rect 14786 14118 14792 14170
rect 14816 14118 14838 14170
rect 14838 14118 14850 14170
rect 14850 14118 14872 14170
rect 14896 14118 14902 14170
rect 14902 14118 14914 14170
rect 14914 14118 14952 14170
rect 14976 14118 14978 14170
rect 14978 14118 15030 14170
rect 15030 14118 15032 14170
rect 14656 14116 14712 14118
rect 14736 14116 14792 14118
rect 14816 14116 14872 14118
rect 14896 14116 14952 14118
rect 14976 14116 15032 14118
rect 13916 13626 13972 13628
rect 13996 13626 14052 13628
rect 14076 13626 14132 13628
rect 14156 13626 14212 13628
rect 14236 13626 14292 13628
rect 13916 13574 13918 13626
rect 13918 13574 13970 13626
rect 13970 13574 13972 13626
rect 13996 13574 14034 13626
rect 14034 13574 14046 13626
rect 14046 13574 14052 13626
rect 14076 13574 14098 13626
rect 14098 13574 14110 13626
rect 14110 13574 14132 13626
rect 14156 13574 14162 13626
rect 14162 13574 14174 13626
rect 14174 13574 14212 13626
rect 14236 13574 14238 13626
rect 14238 13574 14290 13626
rect 14290 13574 14292 13626
rect 13916 13572 13972 13574
rect 13996 13572 14052 13574
rect 14076 13572 14132 13574
rect 14156 13572 14212 13574
rect 14236 13572 14292 13574
rect 14278 12844 14334 12880
rect 14278 12824 14280 12844
rect 14280 12824 14332 12844
rect 14332 12824 14334 12844
rect 13916 12538 13972 12540
rect 13996 12538 14052 12540
rect 14076 12538 14132 12540
rect 14156 12538 14212 12540
rect 14236 12538 14292 12540
rect 13916 12486 13918 12538
rect 13918 12486 13970 12538
rect 13970 12486 13972 12538
rect 13996 12486 14034 12538
rect 14034 12486 14046 12538
rect 14046 12486 14052 12538
rect 14076 12486 14098 12538
rect 14098 12486 14110 12538
rect 14110 12486 14132 12538
rect 14156 12486 14162 12538
rect 14162 12486 14174 12538
rect 14174 12486 14212 12538
rect 14236 12486 14238 12538
rect 14238 12486 14290 12538
rect 14290 12486 14292 12538
rect 13916 12484 13972 12486
rect 13996 12484 14052 12486
rect 14076 12484 14132 12486
rect 14156 12484 14212 12486
rect 14236 12484 14292 12486
rect 12438 7656 12494 7712
rect 11334 3984 11390 4040
rect 11610 3476 11612 3496
rect 11612 3476 11664 3496
rect 11664 3476 11666 3496
rect 11610 3440 11666 3476
rect 13450 6704 13506 6760
rect 13916 11450 13972 11452
rect 13996 11450 14052 11452
rect 14076 11450 14132 11452
rect 14156 11450 14212 11452
rect 14236 11450 14292 11452
rect 13916 11398 13918 11450
rect 13918 11398 13970 11450
rect 13970 11398 13972 11450
rect 13996 11398 14034 11450
rect 14034 11398 14046 11450
rect 14046 11398 14052 11450
rect 14076 11398 14098 11450
rect 14098 11398 14110 11450
rect 14110 11398 14132 11450
rect 14156 11398 14162 11450
rect 14162 11398 14174 11450
rect 14174 11398 14212 11450
rect 14236 11398 14238 11450
rect 14238 11398 14290 11450
rect 14290 11398 14292 11450
rect 13916 11396 13972 11398
rect 13996 11396 14052 11398
rect 14076 11396 14132 11398
rect 14156 11396 14212 11398
rect 14236 11396 14292 11398
rect 13916 10362 13972 10364
rect 13996 10362 14052 10364
rect 14076 10362 14132 10364
rect 14156 10362 14212 10364
rect 14236 10362 14292 10364
rect 13916 10310 13918 10362
rect 13918 10310 13970 10362
rect 13970 10310 13972 10362
rect 13996 10310 14034 10362
rect 14034 10310 14046 10362
rect 14046 10310 14052 10362
rect 14076 10310 14098 10362
rect 14098 10310 14110 10362
rect 14110 10310 14132 10362
rect 14156 10310 14162 10362
rect 14162 10310 14174 10362
rect 14174 10310 14212 10362
rect 14236 10310 14238 10362
rect 14238 10310 14290 10362
rect 14290 10310 14292 10362
rect 13916 10308 13972 10310
rect 13996 10308 14052 10310
rect 14076 10308 14132 10310
rect 14156 10308 14212 10310
rect 14236 10308 14292 10310
rect 14278 10104 14334 10160
rect 14186 9596 14188 9616
rect 14188 9596 14240 9616
rect 14240 9596 14242 9616
rect 14186 9560 14242 9596
rect 14278 9424 14334 9480
rect 14656 13082 14712 13084
rect 14736 13082 14792 13084
rect 14816 13082 14872 13084
rect 14896 13082 14952 13084
rect 14976 13082 15032 13084
rect 14656 13030 14658 13082
rect 14658 13030 14710 13082
rect 14710 13030 14712 13082
rect 14736 13030 14774 13082
rect 14774 13030 14786 13082
rect 14786 13030 14792 13082
rect 14816 13030 14838 13082
rect 14838 13030 14850 13082
rect 14850 13030 14872 13082
rect 14896 13030 14902 13082
rect 14902 13030 14914 13082
rect 14914 13030 14952 13082
rect 14976 13030 14978 13082
rect 14978 13030 15030 13082
rect 15030 13030 15032 13082
rect 14656 13028 14712 13030
rect 14736 13028 14792 13030
rect 14816 13028 14872 13030
rect 14896 13028 14952 13030
rect 14976 13028 15032 13030
rect 14656 11994 14712 11996
rect 14736 11994 14792 11996
rect 14816 11994 14872 11996
rect 14896 11994 14952 11996
rect 14976 11994 15032 11996
rect 14656 11942 14658 11994
rect 14658 11942 14710 11994
rect 14710 11942 14712 11994
rect 14736 11942 14774 11994
rect 14774 11942 14786 11994
rect 14786 11942 14792 11994
rect 14816 11942 14838 11994
rect 14838 11942 14850 11994
rect 14850 11942 14872 11994
rect 14896 11942 14902 11994
rect 14902 11942 14914 11994
rect 14914 11942 14952 11994
rect 14976 11942 14978 11994
rect 14978 11942 15030 11994
rect 15030 11942 15032 11994
rect 14656 11940 14712 11942
rect 14736 11940 14792 11942
rect 14816 11940 14872 11942
rect 14896 11940 14952 11942
rect 14976 11940 15032 11942
rect 16026 14864 16082 14920
rect 15566 12844 15622 12880
rect 15566 12824 15568 12844
rect 15568 12824 15620 12844
rect 15620 12824 15622 12844
rect 14462 10240 14518 10296
rect 14656 10906 14712 10908
rect 14736 10906 14792 10908
rect 14816 10906 14872 10908
rect 14896 10906 14952 10908
rect 14976 10906 15032 10908
rect 14656 10854 14658 10906
rect 14658 10854 14710 10906
rect 14710 10854 14712 10906
rect 14736 10854 14774 10906
rect 14774 10854 14786 10906
rect 14786 10854 14792 10906
rect 14816 10854 14838 10906
rect 14838 10854 14850 10906
rect 14850 10854 14872 10906
rect 14896 10854 14902 10906
rect 14902 10854 14914 10906
rect 14914 10854 14952 10906
rect 14976 10854 14978 10906
rect 14978 10854 15030 10906
rect 15030 10854 15032 10906
rect 14656 10852 14712 10854
rect 14736 10852 14792 10854
rect 14816 10852 14872 10854
rect 14896 10852 14952 10854
rect 14976 10852 15032 10854
rect 14656 9818 14712 9820
rect 14736 9818 14792 9820
rect 14816 9818 14872 9820
rect 14896 9818 14952 9820
rect 14976 9818 15032 9820
rect 14656 9766 14658 9818
rect 14658 9766 14710 9818
rect 14710 9766 14712 9818
rect 14736 9766 14774 9818
rect 14774 9766 14786 9818
rect 14786 9766 14792 9818
rect 14816 9766 14838 9818
rect 14838 9766 14850 9818
rect 14850 9766 14872 9818
rect 14896 9766 14902 9818
rect 14902 9766 14914 9818
rect 14914 9766 14952 9818
rect 14976 9766 14978 9818
rect 14978 9766 15030 9818
rect 15030 9766 15032 9818
rect 14656 9764 14712 9766
rect 14736 9764 14792 9766
rect 14816 9764 14872 9766
rect 14896 9764 14952 9766
rect 14976 9764 15032 9766
rect 13916 9274 13972 9276
rect 13996 9274 14052 9276
rect 14076 9274 14132 9276
rect 14156 9274 14212 9276
rect 14236 9274 14292 9276
rect 13916 9222 13918 9274
rect 13918 9222 13970 9274
rect 13970 9222 13972 9274
rect 13996 9222 14034 9274
rect 14034 9222 14046 9274
rect 14046 9222 14052 9274
rect 14076 9222 14098 9274
rect 14098 9222 14110 9274
rect 14110 9222 14132 9274
rect 14156 9222 14162 9274
rect 14162 9222 14174 9274
rect 14174 9222 14212 9274
rect 14236 9222 14238 9274
rect 14238 9222 14290 9274
rect 14290 9222 14292 9274
rect 13916 9220 13972 9222
rect 13996 9220 14052 9222
rect 14076 9220 14132 9222
rect 14156 9220 14212 9222
rect 14236 9220 14292 9222
rect 15750 9580 15806 9616
rect 15750 9560 15752 9580
rect 15752 9560 15804 9580
rect 15804 9560 15806 9580
rect 14656 8730 14712 8732
rect 14736 8730 14792 8732
rect 14816 8730 14872 8732
rect 14896 8730 14952 8732
rect 14976 8730 15032 8732
rect 14656 8678 14658 8730
rect 14658 8678 14710 8730
rect 14710 8678 14712 8730
rect 14736 8678 14774 8730
rect 14774 8678 14786 8730
rect 14786 8678 14792 8730
rect 14816 8678 14838 8730
rect 14838 8678 14850 8730
rect 14850 8678 14872 8730
rect 14896 8678 14902 8730
rect 14902 8678 14914 8730
rect 14914 8678 14952 8730
rect 14976 8678 14978 8730
rect 14978 8678 15030 8730
rect 15030 8678 15032 8730
rect 14656 8676 14712 8678
rect 14736 8676 14792 8678
rect 14816 8676 14872 8678
rect 14896 8676 14952 8678
rect 14976 8676 15032 8678
rect 13916 8186 13972 8188
rect 13996 8186 14052 8188
rect 14076 8186 14132 8188
rect 14156 8186 14212 8188
rect 14236 8186 14292 8188
rect 13916 8134 13918 8186
rect 13918 8134 13970 8186
rect 13970 8134 13972 8186
rect 13996 8134 14034 8186
rect 14034 8134 14046 8186
rect 14046 8134 14052 8186
rect 14076 8134 14098 8186
rect 14098 8134 14110 8186
rect 14110 8134 14132 8186
rect 14156 8134 14162 8186
rect 14162 8134 14174 8186
rect 14174 8134 14212 8186
rect 14236 8134 14238 8186
rect 14238 8134 14290 8186
rect 14290 8134 14292 8186
rect 13916 8132 13972 8134
rect 13996 8132 14052 8134
rect 14076 8132 14132 8134
rect 14156 8132 14212 8134
rect 14236 8132 14292 8134
rect 13916 7098 13972 7100
rect 13996 7098 14052 7100
rect 14076 7098 14132 7100
rect 14156 7098 14212 7100
rect 14236 7098 14292 7100
rect 13916 7046 13918 7098
rect 13918 7046 13970 7098
rect 13970 7046 13972 7098
rect 13996 7046 14034 7098
rect 14034 7046 14046 7098
rect 14046 7046 14052 7098
rect 14076 7046 14098 7098
rect 14098 7046 14110 7098
rect 14110 7046 14132 7098
rect 14156 7046 14162 7098
rect 14162 7046 14174 7098
rect 14174 7046 14212 7098
rect 14236 7046 14238 7098
rect 14238 7046 14290 7098
rect 14290 7046 14292 7098
rect 13916 7044 13972 7046
rect 13996 7044 14052 7046
rect 14076 7044 14132 7046
rect 14156 7044 14212 7046
rect 14236 7044 14292 7046
rect 14370 6860 14426 6896
rect 14370 6840 14372 6860
rect 14372 6840 14424 6860
rect 14424 6840 14426 6860
rect 14656 7642 14712 7644
rect 14736 7642 14792 7644
rect 14816 7642 14872 7644
rect 14896 7642 14952 7644
rect 14976 7642 15032 7644
rect 14656 7590 14658 7642
rect 14658 7590 14710 7642
rect 14710 7590 14712 7642
rect 14736 7590 14774 7642
rect 14774 7590 14786 7642
rect 14786 7590 14792 7642
rect 14816 7590 14838 7642
rect 14838 7590 14850 7642
rect 14850 7590 14872 7642
rect 14896 7590 14902 7642
rect 14902 7590 14914 7642
rect 14914 7590 14952 7642
rect 14976 7590 14978 7642
rect 14978 7590 15030 7642
rect 15030 7590 15032 7642
rect 14656 7588 14712 7590
rect 14736 7588 14792 7590
rect 14816 7588 14872 7590
rect 14896 7588 14952 7590
rect 14976 7588 15032 7590
rect 14002 6740 14004 6760
rect 14004 6740 14056 6760
rect 14056 6740 14058 6760
rect 14002 6704 14058 6740
rect 15566 6704 15622 6760
rect 14656 6554 14712 6556
rect 14736 6554 14792 6556
rect 14816 6554 14872 6556
rect 14896 6554 14952 6556
rect 14976 6554 15032 6556
rect 14656 6502 14658 6554
rect 14658 6502 14710 6554
rect 14710 6502 14712 6554
rect 14736 6502 14774 6554
rect 14774 6502 14786 6554
rect 14786 6502 14792 6554
rect 14816 6502 14838 6554
rect 14838 6502 14850 6554
rect 14850 6502 14872 6554
rect 14896 6502 14902 6554
rect 14902 6502 14914 6554
rect 14914 6502 14952 6554
rect 14976 6502 14978 6554
rect 14978 6502 15030 6554
rect 15030 6502 15032 6554
rect 14656 6500 14712 6502
rect 14736 6500 14792 6502
rect 14816 6500 14872 6502
rect 14896 6500 14952 6502
rect 14976 6500 15032 6502
rect 14462 6432 14518 6488
rect 13916 6010 13972 6012
rect 13996 6010 14052 6012
rect 14076 6010 14132 6012
rect 14156 6010 14212 6012
rect 14236 6010 14292 6012
rect 13916 5958 13918 6010
rect 13918 5958 13970 6010
rect 13970 5958 13972 6010
rect 13996 5958 14034 6010
rect 14034 5958 14046 6010
rect 14046 5958 14052 6010
rect 14076 5958 14098 6010
rect 14098 5958 14110 6010
rect 14110 5958 14132 6010
rect 14156 5958 14162 6010
rect 14162 5958 14174 6010
rect 14174 5958 14212 6010
rect 14236 5958 14238 6010
rect 14238 5958 14290 6010
rect 14290 5958 14292 6010
rect 13916 5956 13972 5958
rect 13996 5956 14052 5958
rect 14076 5956 14132 5958
rect 14156 5956 14212 5958
rect 14236 5956 14292 5958
rect 13916 4922 13972 4924
rect 13996 4922 14052 4924
rect 14076 4922 14132 4924
rect 14156 4922 14212 4924
rect 14236 4922 14292 4924
rect 13916 4870 13918 4922
rect 13918 4870 13970 4922
rect 13970 4870 13972 4922
rect 13996 4870 14034 4922
rect 14034 4870 14046 4922
rect 14046 4870 14052 4922
rect 14076 4870 14098 4922
rect 14098 4870 14110 4922
rect 14110 4870 14132 4922
rect 14156 4870 14162 4922
rect 14162 4870 14174 4922
rect 14174 4870 14212 4922
rect 14236 4870 14238 4922
rect 14238 4870 14290 4922
rect 14290 4870 14292 4922
rect 13916 4868 13972 4870
rect 13996 4868 14052 4870
rect 14076 4868 14132 4870
rect 14156 4868 14212 4870
rect 14236 4868 14292 4870
rect 14656 5466 14712 5468
rect 14736 5466 14792 5468
rect 14816 5466 14872 5468
rect 14896 5466 14952 5468
rect 14976 5466 15032 5468
rect 14656 5414 14658 5466
rect 14658 5414 14710 5466
rect 14710 5414 14712 5466
rect 14736 5414 14774 5466
rect 14774 5414 14786 5466
rect 14786 5414 14792 5466
rect 14816 5414 14838 5466
rect 14838 5414 14850 5466
rect 14850 5414 14872 5466
rect 14896 5414 14902 5466
rect 14902 5414 14914 5466
rect 14914 5414 14952 5466
rect 14976 5414 14978 5466
rect 14978 5414 15030 5466
rect 15030 5414 15032 5466
rect 14656 5412 14712 5414
rect 14736 5412 14792 5414
rect 14816 5412 14872 5414
rect 14896 5412 14952 5414
rect 14976 5412 15032 5414
rect 13916 3834 13972 3836
rect 13996 3834 14052 3836
rect 14076 3834 14132 3836
rect 14156 3834 14212 3836
rect 14236 3834 14292 3836
rect 13916 3782 13918 3834
rect 13918 3782 13970 3834
rect 13970 3782 13972 3834
rect 13996 3782 14034 3834
rect 14034 3782 14046 3834
rect 14046 3782 14052 3834
rect 14076 3782 14098 3834
rect 14098 3782 14110 3834
rect 14110 3782 14132 3834
rect 14156 3782 14162 3834
rect 14162 3782 14174 3834
rect 14174 3782 14212 3834
rect 14236 3782 14238 3834
rect 14238 3782 14290 3834
rect 14290 3782 14292 3834
rect 13916 3780 13972 3782
rect 13996 3780 14052 3782
rect 14076 3780 14132 3782
rect 14156 3780 14212 3782
rect 14236 3780 14292 3782
rect 14656 4378 14712 4380
rect 14736 4378 14792 4380
rect 14816 4378 14872 4380
rect 14896 4378 14952 4380
rect 14976 4378 15032 4380
rect 14656 4326 14658 4378
rect 14658 4326 14710 4378
rect 14710 4326 14712 4378
rect 14736 4326 14774 4378
rect 14774 4326 14786 4378
rect 14786 4326 14792 4378
rect 14816 4326 14838 4378
rect 14838 4326 14850 4378
rect 14850 4326 14872 4378
rect 14896 4326 14902 4378
rect 14902 4326 14914 4378
rect 14914 4326 14952 4378
rect 14976 4326 14978 4378
rect 14978 4326 15030 4378
rect 15030 4326 15032 4378
rect 14656 4324 14712 4326
rect 14736 4324 14792 4326
rect 14816 4324 14872 4326
rect 14896 4324 14952 4326
rect 14976 4324 15032 4326
rect 16578 10376 16634 10432
rect 16486 6296 16542 6352
rect 16670 6160 16726 6216
rect 14656 3290 14712 3292
rect 14736 3290 14792 3292
rect 14816 3290 14872 3292
rect 14896 3290 14952 3292
rect 14976 3290 15032 3292
rect 14656 3238 14658 3290
rect 14658 3238 14710 3290
rect 14710 3238 14712 3290
rect 14736 3238 14774 3290
rect 14774 3238 14786 3290
rect 14786 3238 14792 3290
rect 14816 3238 14838 3290
rect 14838 3238 14850 3290
rect 14850 3238 14872 3290
rect 14896 3238 14902 3290
rect 14902 3238 14914 3290
rect 14914 3238 14952 3290
rect 14976 3238 14978 3290
rect 14978 3238 15030 3290
rect 15030 3238 15032 3290
rect 14656 3236 14712 3238
rect 14736 3236 14792 3238
rect 14816 3236 14872 3238
rect 14896 3236 14952 3238
rect 14976 3236 15032 3238
rect 15750 3440 15806 3496
rect 13916 2746 13972 2748
rect 13996 2746 14052 2748
rect 14076 2746 14132 2748
rect 14156 2746 14212 2748
rect 14236 2746 14292 2748
rect 13916 2694 13918 2746
rect 13918 2694 13970 2746
rect 13970 2694 13972 2746
rect 13996 2694 14034 2746
rect 14034 2694 14046 2746
rect 14046 2694 14052 2746
rect 14076 2694 14098 2746
rect 14098 2694 14110 2746
rect 14110 2694 14132 2746
rect 14156 2694 14162 2746
rect 14162 2694 14174 2746
rect 14174 2694 14212 2746
rect 14236 2694 14238 2746
rect 14238 2694 14290 2746
rect 14290 2694 14292 2746
rect 13916 2692 13972 2694
rect 13996 2692 14052 2694
rect 14076 2692 14132 2694
rect 14156 2692 14212 2694
rect 14236 2692 14292 2694
rect 1398 2216 1454 2272
rect 2656 2202 2712 2204
rect 2736 2202 2792 2204
rect 2816 2202 2872 2204
rect 2896 2202 2952 2204
rect 2976 2202 3032 2204
rect 2656 2150 2658 2202
rect 2658 2150 2710 2202
rect 2710 2150 2712 2202
rect 2736 2150 2774 2202
rect 2774 2150 2786 2202
rect 2786 2150 2792 2202
rect 2816 2150 2838 2202
rect 2838 2150 2850 2202
rect 2850 2150 2872 2202
rect 2896 2150 2902 2202
rect 2902 2150 2914 2202
rect 2914 2150 2952 2202
rect 2976 2150 2978 2202
rect 2978 2150 3030 2202
rect 3030 2150 3032 2202
rect 2656 2148 2712 2150
rect 2736 2148 2792 2150
rect 2816 2148 2872 2150
rect 2896 2148 2952 2150
rect 2976 2148 3032 2150
rect 8656 2202 8712 2204
rect 8736 2202 8792 2204
rect 8816 2202 8872 2204
rect 8896 2202 8952 2204
rect 8976 2202 9032 2204
rect 8656 2150 8658 2202
rect 8658 2150 8710 2202
rect 8710 2150 8712 2202
rect 8736 2150 8774 2202
rect 8774 2150 8786 2202
rect 8786 2150 8792 2202
rect 8816 2150 8838 2202
rect 8838 2150 8850 2202
rect 8850 2150 8872 2202
rect 8896 2150 8902 2202
rect 8902 2150 8914 2202
rect 8914 2150 8952 2202
rect 8976 2150 8978 2202
rect 8978 2150 9030 2202
rect 9030 2150 9032 2202
rect 8656 2148 8712 2150
rect 8736 2148 8792 2150
rect 8816 2148 8872 2150
rect 8896 2148 8952 2150
rect 8976 2148 9032 2150
rect 14656 2202 14712 2204
rect 14736 2202 14792 2204
rect 14816 2202 14872 2204
rect 14896 2202 14952 2204
rect 14976 2202 15032 2204
rect 14656 2150 14658 2202
rect 14658 2150 14710 2202
rect 14710 2150 14712 2202
rect 14736 2150 14774 2202
rect 14774 2150 14786 2202
rect 14786 2150 14792 2202
rect 14816 2150 14838 2202
rect 14838 2150 14850 2202
rect 14850 2150 14872 2202
rect 14896 2150 14902 2202
rect 14902 2150 14914 2202
rect 14914 2150 14952 2202
rect 14976 2150 14978 2202
rect 14978 2150 15030 2202
rect 15030 2150 15032 2202
rect 14656 2148 14712 2150
rect 14736 2148 14792 2150
rect 14816 2148 14872 2150
rect 14896 2148 14952 2150
rect 14976 2148 15032 2150
<< metal3 >>
rect 0 18594 800 18624
rect 1209 18594 1275 18597
rect 0 18592 1275 18594
rect 0 18536 1214 18592
rect 1270 18536 1275 18592
rect 0 18534 1275 18536
rect 0 18504 800 18534
rect 1209 18531 1275 18534
rect 2646 18528 3042 18529
rect 2646 18464 2652 18528
rect 2716 18464 2732 18528
rect 2796 18464 2812 18528
rect 2876 18464 2892 18528
rect 2956 18464 2972 18528
rect 3036 18464 3042 18528
rect 2646 18463 3042 18464
rect 8646 18528 9042 18529
rect 8646 18464 8652 18528
rect 8716 18464 8732 18528
rect 8796 18464 8812 18528
rect 8876 18464 8892 18528
rect 8956 18464 8972 18528
rect 9036 18464 9042 18528
rect 8646 18463 9042 18464
rect 14646 18528 15042 18529
rect 14646 18464 14652 18528
rect 14716 18464 14732 18528
rect 14796 18464 14812 18528
rect 14876 18464 14892 18528
rect 14956 18464 14972 18528
rect 15036 18464 15042 18528
rect 14646 18463 15042 18464
rect 12433 18050 12499 18053
rect 12566 18050 12572 18052
rect 12433 18048 12572 18050
rect 12433 17992 12438 18048
rect 12494 17992 12572 18048
rect 12433 17990 12572 17992
rect 12433 17987 12499 17990
rect 12566 17988 12572 17990
rect 12636 17988 12642 18052
rect 1906 17984 2302 17985
rect 1906 17920 1912 17984
rect 1976 17920 1992 17984
rect 2056 17920 2072 17984
rect 2136 17920 2152 17984
rect 2216 17920 2232 17984
rect 2296 17920 2302 17984
rect 1906 17919 2302 17920
rect 7906 17984 8302 17985
rect 7906 17920 7912 17984
rect 7976 17920 7992 17984
rect 8056 17920 8072 17984
rect 8136 17920 8152 17984
rect 8216 17920 8232 17984
rect 8296 17920 8302 17984
rect 7906 17919 8302 17920
rect 13906 17984 14302 17985
rect 13906 17920 13912 17984
rect 13976 17920 13992 17984
rect 14056 17920 14072 17984
rect 14136 17920 14152 17984
rect 14216 17920 14232 17984
rect 14296 17920 14302 17984
rect 13906 17919 14302 17920
rect 0 17506 800 17536
rect 1301 17506 1367 17509
rect 0 17504 1367 17506
rect 0 17448 1306 17504
rect 1362 17448 1367 17504
rect 0 17446 1367 17448
rect 0 17416 800 17446
rect 1301 17443 1367 17446
rect 2646 17440 3042 17441
rect 2646 17376 2652 17440
rect 2716 17376 2732 17440
rect 2796 17376 2812 17440
rect 2876 17376 2892 17440
rect 2956 17376 2972 17440
rect 3036 17376 3042 17440
rect 2646 17375 3042 17376
rect 8646 17440 9042 17441
rect 8646 17376 8652 17440
rect 8716 17376 8732 17440
rect 8796 17376 8812 17440
rect 8876 17376 8892 17440
rect 8956 17376 8972 17440
rect 9036 17376 9042 17440
rect 8646 17375 9042 17376
rect 14646 17440 15042 17441
rect 14646 17376 14652 17440
rect 14716 17376 14732 17440
rect 14796 17376 14812 17440
rect 14876 17376 14892 17440
rect 14956 17376 14972 17440
rect 15036 17376 15042 17440
rect 14646 17375 15042 17376
rect 1906 16896 2302 16897
rect 1906 16832 1912 16896
rect 1976 16832 1992 16896
rect 2056 16832 2072 16896
rect 2136 16832 2152 16896
rect 2216 16832 2232 16896
rect 2296 16832 2302 16896
rect 1906 16831 2302 16832
rect 7906 16896 8302 16897
rect 7906 16832 7912 16896
rect 7976 16832 7992 16896
rect 8056 16832 8072 16896
rect 8136 16832 8152 16896
rect 8216 16832 8232 16896
rect 8296 16832 8302 16896
rect 7906 16831 8302 16832
rect 13906 16896 14302 16897
rect 13906 16832 13912 16896
rect 13976 16832 13992 16896
rect 14056 16832 14072 16896
rect 14136 16832 14152 16896
rect 14216 16832 14232 16896
rect 14296 16832 14302 16896
rect 13906 16831 14302 16832
rect 841 16554 907 16557
rect 798 16552 907 16554
rect 798 16496 846 16552
rect 902 16496 907 16552
rect 798 16491 907 16496
rect 798 16448 858 16491
rect 0 16358 858 16448
rect 0 16328 800 16358
rect 2646 16352 3042 16353
rect 2646 16288 2652 16352
rect 2716 16288 2732 16352
rect 2796 16288 2812 16352
rect 2876 16288 2892 16352
rect 2956 16288 2972 16352
rect 3036 16288 3042 16352
rect 2646 16287 3042 16288
rect 8646 16352 9042 16353
rect 8646 16288 8652 16352
rect 8716 16288 8732 16352
rect 8796 16288 8812 16352
rect 8876 16288 8892 16352
rect 8956 16288 8972 16352
rect 9036 16288 9042 16352
rect 8646 16287 9042 16288
rect 14646 16352 15042 16353
rect 14646 16288 14652 16352
rect 14716 16288 14732 16352
rect 14796 16288 14812 16352
rect 14876 16288 14892 16352
rect 14956 16288 14972 16352
rect 15036 16288 15042 16352
rect 14646 16287 15042 16288
rect 1906 15808 2302 15809
rect 1906 15744 1912 15808
rect 1976 15744 1992 15808
rect 2056 15744 2072 15808
rect 2136 15744 2152 15808
rect 2216 15744 2232 15808
rect 2296 15744 2302 15808
rect 1906 15743 2302 15744
rect 7906 15808 8302 15809
rect 7906 15744 7912 15808
rect 7976 15744 7992 15808
rect 8056 15744 8072 15808
rect 8136 15744 8152 15808
rect 8216 15744 8232 15808
rect 8296 15744 8302 15808
rect 7906 15743 8302 15744
rect 13906 15808 14302 15809
rect 13906 15744 13912 15808
rect 13976 15744 13992 15808
rect 14056 15744 14072 15808
rect 14136 15744 14152 15808
rect 14216 15744 14232 15808
rect 14296 15744 14302 15808
rect 13906 15743 14302 15744
rect 12065 15602 12131 15605
rect 12709 15602 12775 15605
rect 12065 15600 12775 15602
rect 12065 15544 12070 15600
rect 12126 15544 12714 15600
rect 12770 15544 12775 15600
rect 12065 15542 12775 15544
rect 12065 15539 12131 15542
rect 12709 15539 12775 15542
rect 841 15466 907 15469
rect 798 15464 907 15466
rect 798 15408 846 15464
rect 902 15408 907 15464
rect 798 15403 907 15408
rect 798 15360 858 15403
rect 0 15270 858 15360
rect 0 15240 800 15270
rect 2646 15264 3042 15265
rect 2646 15200 2652 15264
rect 2716 15200 2732 15264
rect 2796 15200 2812 15264
rect 2876 15200 2892 15264
rect 2956 15200 2972 15264
rect 3036 15200 3042 15264
rect 2646 15199 3042 15200
rect 8646 15264 9042 15265
rect 8646 15200 8652 15264
rect 8716 15200 8732 15264
rect 8796 15200 8812 15264
rect 8876 15200 8892 15264
rect 8956 15200 8972 15264
rect 9036 15200 9042 15264
rect 8646 15199 9042 15200
rect 14646 15264 15042 15265
rect 14646 15200 14652 15264
rect 14716 15200 14732 15264
rect 14796 15200 14812 15264
rect 14876 15200 14892 15264
rect 14956 15200 14972 15264
rect 15036 15200 15042 15264
rect 14646 15199 15042 15200
rect 3233 14922 3299 14925
rect 16021 14922 16087 14925
rect 3233 14920 16087 14922
rect 3233 14864 3238 14920
rect 3294 14864 16026 14920
rect 16082 14864 16087 14920
rect 3233 14862 16087 14864
rect 3233 14859 3299 14862
rect 16021 14859 16087 14862
rect 1906 14720 2302 14721
rect 1906 14656 1912 14720
rect 1976 14656 1992 14720
rect 2056 14656 2072 14720
rect 2136 14656 2152 14720
rect 2216 14656 2232 14720
rect 2296 14656 2302 14720
rect 1906 14655 2302 14656
rect 7906 14720 8302 14721
rect 7906 14656 7912 14720
rect 7976 14656 7992 14720
rect 8056 14656 8072 14720
rect 8136 14656 8152 14720
rect 8216 14656 8232 14720
rect 8296 14656 8302 14720
rect 7906 14655 8302 14656
rect 13906 14720 14302 14721
rect 13906 14656 13912 14720
rect 13976 14656 13992 14720
rect 14056 14656 14072 14720
rect 14136 14656 14152 14720
rect 14216 14656 14232 14720
rect 14296 14656 14302 14720
rect 13906 14655 14302 14656
rect 841 14378 907 14381
rect 798 14376 907 14378
rect 798 14320 846 14376
rect 902 14320 907 14376
rect 798 14315 907 14320
rect 798 14272 858 14315
rect 0 14182 858 14272
rect 0 14152 800 14182
rect 2646 14176 3042 14177
rect 2646 14112 2652 14176
rect 2716 14112 2732 14176
rect 2796 14112 2812 14176
rect 2876 14112 2892 14176
rect 2956 14112 2972 14176
rect 3036 14112 3042 14176
rect 2646 14111 3042 14112
rect 8646 14176 9042 14177
rect 8646 14112 8652 14176
rect 8716 14112 8732 14176
rect 8796 14112 8812 14176
rect 8876 14112 8892 14176
rect 8956 14112 8972 14176
rect 9036 14112 9042 14176
rect 8646 14111 9042 14112
rect 14646 14176 15042 14177
rect 14646 14112 14652 14176
rect 14716 14112 14732 14176
rect 14796 14112 14812 14176
rect 14876 14112 14892 14176
rect 14956 14112 14972 14176
rect 15036 14112 15042 14176
rect 14646 14111 15042 14112
rect 1906 13632 2302 13633
rect 1906 13568 1912 13632
rect 1976 13568 1992 13632
rect 2056 13568 2072 13632
rect 2136 13568 2152 13632
rect 2216 13568 2232 13632
rect 2296 13568 2302 13632
rect 1906 13567 2302 13568
rect 7906 13632 8302 13633
rect 7906 13568 7912 13632
rect 7976 13568 7992 13632
rect 8056 13568 8072 13632
rect 8136 13568 8152 13632
rect 8216 13568 8232 13632
rect 8296 13568 8302 13632
rect 7906 13567 8302 13568
rect 13906 13632 14302 13633
rect 13906 13568 13912 13632
rect 13976 13568 13992 13632
rect 14056 13568 14072 13632
rect 14136 13568 14152 13632
rect 14216 13568 14232 13632
rect 14296 13568 14302 13632
rect 13906 13567 14302 13568
rect 841 13290 907 13293
rect 798 13288 907 13290
rect 798 13232 846 13288
rect 902 13232 907 13288
rect 798 13227 907 13232
rect 798 13184 858 13227
rect 0 13094 858 13184
rect 0 13064 800 13094
rect 2646 13088 3042 13089
rect 2646 13024 2652 13088
rect 2716 13024 2732 13088
rect 2796 13024 2812 13088
rect 2876 13024 2892 13088
rect 2956 13024 2972 13088
rect 3036 13024 3042 13088
rect 2646 13023 3042 13024
rect 8646 13088 9042 13089
rect 8646 13024 8652 13088
rect 8716 13024 8732 13088
rect 8796 13024 8812 13088
rect 8876 13024 8892 13088
rect 8956 13024 8972 13088
rect 9036 13024 9042 13088
rect 8646 13023 9042 13024
rect 14646 13088 15042 13089
rect 14646 13024 14652 13088
rect 14716 13024 14732 13088
rect 14796 13024 14812 13088
rect 14876 13024 14892 13088
rect 14956 13024 14972 13088
rect 15036 13024 15042 13088
rect 14646 13023 15042 13024
rect 14273 12882 14339 12885
rect 15561 12882 15627 12885
rect 14273 12880 15627 12882
rect 14273 12824 14278 12880
rect 14334 12824 15566 12880
rect 15622 12824 15627 12880
rect 14273 12822 15627 12824
rect 14273 12819 14339 12822
rect 15561 12819 15627 12822
rect 1906 12544 2302 12545
rect 1906 12480 1912 12544
rect 1976 12480 1992 12544
rect 2056 12480 2072 12544
rect 2136 12480 2152 12544
rect 2216 12480 2232 12544
rect 2296 12480 2302 12544
rect 1906 12479 2302 12480
rect 7906 12544 8302 12545
rect 7906 12480 7912 12544
rect 7976 12480 7992 12544
rect 8056 12480 8072 12544
rect 8136 12480 8152 12544
rect 8216 12480 8232 12544
rect 8296 12480 8302 12544
rect 7906 12479 8302 12480
rect 13906 12544 14302 12545
rect 13906 12480 13912 12544
rect 13976 12480 13992 12544
rect 14056 12480 14072 12544
rect 14136 12480 14152 12544
rect 14216 12480 14232 12544
rect 14296 12480 14302 12544
rect 13906 12479 14302 12480
rect 841 12202 907 12205
rect 798 12200 907 12202
rect 798 12144 846 12200
rect 902 12144 907 12200
rect 798 12139 907 12144
rect 798 12096 858 12139
rect 0 12006 858 12096
rect 0 11976 800 12006
rect 2646 12000 3042 12001
rect 2646 11936 2652 12000
rect 2716 11936 2732 12000
rect 2796 11936 2812 12000
rect 2876 11936 2892 12000
rect 2956 11936 2972 12000
rect 3036 11936 3042 12000
rect 2646 11935 3042 11936
rect 8646 12000 9042 12001
rect 8646 11936 8652 12000
rect 8716 11936 8732 12000
rect 8796 11936 8812 12000
rect 8876 11936 8892 12000
rect 8956 11936 8972 12000
rect 9036 11936 9042 12000
rect 8646 11935 9042 11936
rect 14646 12000 15042 12001
rect 14646 11936 14652 12000
rect 14716 11936 14732 12000
rect 14796 11936 14812 12000
rect 14876 11936 14892 12000
rect 14956 11936 14972 12000
rect 15036 11936 15042 12000
rect 14646 11935 15042 11936
rect 1906 11456 2302 11457
rect 1906 11392 1912 11456
rect 1976 11392 1992 11456
rect 2056 11392 2072 11456
rect 2136 11392 2152 11456
rect 2216 11392 2232 11456
rect 2296 11392 2302 11456
rect 1906 11391 2302 11392
rect 7906 11456 8302 11457
rect 7906 11392 7912 11456
rect 7976 11392 7992 11456
rect 8056 11392 8072 11456
rect 8136 11392 8152 11456
rect 8216 11392 8232 11456
rect 8296 11392 8302 11456
rect 7906 11391 8302 11392
rect 13906 11456 14302 11457
rect 13906 11392 13912 11456
rect 13976 11392 13992 11456
rect 14056 11392 14072 11456
rect 14136 11392 14152 11456
rect 14216 11392 14232 11456
rect 14296 11392 14302 11456
rect 13906 11391 14302 11392
rect 0 10978 800 11008
rect 1301 10978 1367 10981
rect 0 10976 1367 10978
rect 0 10920 1306 10976
rect 1362 10920 1367 10976
rect 0 10918 1367 10920
rect 0 10888 800 10918
rect 1301 10915 1367 10918
rect 2646 10912 3042 10913
rect 2646 10848 2652 10912
rect 2716 10848 2732 10912
rect 2796 10848 2812 10912
rect 2876 10848 2892 10912
rect 2956 10848 2972 10912
rect 3036 10848 3042 10912
rect 2646 10847 3042 10848
rect 8646 10912 9042 10913
rect 8646 10848 8652 10912
rect 8716 10848 8732 10912
rect 8796 10848 8812 10912
rect 8876 10848 8892 10912
rect 8956 10848 8972 10912
rect 9036 10848 9042 10912
rect 8646 10847 9042 10848
rect 14646 10912 15042 10913
rect 14646 10848 14652 10912
rect 14716 10848 14732 10912
rect 14796 10848 14812 10912
rect 14876 10848 14892 10912
rect 14956 10848 14972 10912
rect 15036 10848 15042 10912
rect 14646 10847 15042 10848
rect 16573 10434 16639 10437
rect 18157 10434 18957 10464
rect 16573 10432 18957 10434
rect 16573 10376 16578 10432
rect 16634 10376 18957 10432
rect 16573 10374 18957 10376
rect 16573 10371 16639 10374
rect 1906 10368 2302 10369
rect 1906 10304 1912 10368
rect 1976 10304 1992 10368
rect 2056 10304 2072 10368
rect 2136 10304 2152 10368
rect 2216 10304 2232 10368
rect 2296 10304 2302 10368
rect 1906 10303 2302 10304
rect 7906 10368 8302 10369
rect 7906 10304 7912 10368
rect 7976 10304 7992 10368
rect 8056 10304 8072 10368
rect 8136 10304 8152 10368
rect 8216 10304 8232 10368
rect 8296 10304 8302 10368
rect 7906 10303 8302 10304
rect 13906 10368 14302 10369
rect 13906 10304 13912 10368
rect 13976 10304 13992 10368
rect 14056 10304 14072 10368
rect 14136 10304 14152 10368
rect 14216 10304 14232 10368
rect 14296 10304 14302 10368
rect 18157 10344 18957 10374
rect 13906 10303 14302 10304
rect 14457 10298 14523 10301
rect 14414 10296 14523 10298
rect 14414 10240 14462 10296
rect 14518 10240 14523 10296
rect 14414 10235 14523 10240
rect 14273 10162 14339 10165
rect 14414 10162 14474 10235
rect 14273 10160 14474 10162
rect 14273 10104 14278 10160
rect 14334 10104 14474 10160
rect 14273 10102 14474 10104
rect 14273 10099 14339 10102
rect 0 9890 800 9920
rect 1301 9890 1367 9893
rect 0 9888 1367 9890
rect 0 9832 1306 9888
rect 1362 9832 1367 9888
rect 0 9830 1367 9832
rect 0 9800 800 9830
rect 1301 9827 1367 9830
rect 2646 9824 3042 9825
rect 2646 9760 2652 9824
rect 2716 9760 2732 9824
rect 2796 9760 2812 9824
rect 2876 9760 2892 9824
rect 2956 9760 2972 9824
rect 3036 9760 3042 9824
rect 2646 9759 3042 9760
rect 8646 9824 9042 9825
rect 8646 9760 8652 9824
rect 8716 9760 8732 9824
rect 8796 9760 8812 9824
rect 8876 9760 8892 9824
rect 8956 9760 8972 9824
rect 9036 9760 9042 9824
rect 8646 9759 9042 9760
rect 14646 9824 15042 9825
rect 14646 9760 14652 9824
rect 14716 9760 14732 9824
rect 14796 9760 14812 9824
rect 14876 9760 14892 9824
rect 14956 9760 14972 9824
rect 15036 9760 15042 9824
rect 14646 9759 15042 9760
rect 14181 9618 14247 9621
rect 15745 9618 15811 9621
rect 14181 9616 15811 9618
rect 14181 9560 14186 9616
rect 14242 9560 15750 9616
rect 15806 9560 15811 9616
rect 14181 9558 15811 9560
rect 14181 9555 14247 9558
rect 15745 9555 15811 9558
rect 14273 9482 14339 9485
rect 14406 9482 14412 9484
rect 14273 9480 14412 9482
rect 14273 9424 14278 9480
rect 14334 9424 14412 9480
rect 14273 9422 14412 9424
rect 14273 9419 14339 9422
rect 14406 9420 14412 9422
rect 14476 9420 14482 9484
rect 1906 9280 2302 9281
rect 1906 9216 1912 9280
rect 1976 9216 1992 9280
rect 2056 9216 2072 9280
rect 2136 9216 2152 9280
rect 2216 9216 2232 9280
rect 2296 9216 2302 9280
rect 1906 9215 2302 9216
rect 7906 9280 8302 9281
rect 7906 9216 7912 9280
rect 7976 9216 7992 9280
rect 8056 9216 8072 9280
rect 8136 9216 8152 9280
rect 8216 9216 8232 9280
rect 8296 9216 8302 9280
rect 7906 9215 8302 9216
rect 13906 9280 14302 9281
rect 13906 9216 13912 9280
rect 13976 9216 13992 9280
rect 14056 9216 14072 9280
rect 14136 9216 14152 9280
rect 14216 9216 14232 9280
rect 14296 9216 14302 9280
rect 13906 9215 14302 9216
rect 0 8802 800 8832
rect 1301 8802 1367 8805
rect 0 8800 1367 8802
rect 0 8744 1306 8800
rect 1362 8744 1367 8800
rect 0 8742 1367 8744
rect 0 8712 800 8742
rect 1301 8739 1367 8742
rect 2646 8736 3042 8737
rect 2646 8672 2652 8736
rect 2716 8672 2732 8736
rect 2796 8672 2812 8736
rect 2876 8672 2892 8736
rect 2956 8672 2972 8736
rect 3036 8672 3042 8736
rect 2646 8671 3042 8672
rect 8646 8736 9042 8737
rect 8646 8672 8652 8736
rect 8716 8672 8732 8736
rect 8796 8672 8812 8736
rect 8876 8672 8892 8736
rect 8956 8672 8972 8736
rect 9036 8672 9042 8736
rect 8646 8671 9042 8672
rect 14646 8736 15042 8737
rect 14646 8672 14652 8736
rect 14716 8672 14732 8736
rect 14796 8672 14812 8736
rect 14876 8672 14892 8736
rect 14956 8672 14972 8736
rect 15036 8672 15042 8736
rect 14646 8671 15042 8672
rect 1906 8192 2302 8193
rect 1906 8128 1912 8192
rect 1976 8128 1992 8192
rect 2056 8128 2072 8192
rect 2136 8128 2152 8192
rect 2216 8128 2232 8192
rect 2296 8128 2302 8192
rect 1906 8127 2302 8128
rect 7906 8192 8302 8193
rect 7906 8128 7912 8192
rect 7976 8128 7992 8192
rect 8056 8128 8072 8192
rect 8136 8128 8152 8192
rect 8216 8128 8232 8192
rect 8296 8128 8302 8192
rect 7906 8127 8302 8128
rect 13906 8192 14302 8193
rect 13906 8128 13912 8192
rect 13976 8128 13992 8192
rect 14056 8128 14072 8192
rect 14136 8128 14152 8192
rect 14216 8128 14232 8192
rect 14296 8128 14302 8192
rect 13906 8127 14302 8128
rect 0 7714 800 7744
rect 1301 7714 1367 7717
rect 0 7712 1367 7714
rect 0 7656 1306 7712
rect 1362 7656 1367 7712
rect 0 7654 1367 7656
rect 0 7624 800 7654
rect 1301 7651 1367 7654
rect 12433 7714 12499 7717
rect 12566 7714 12572 7716
rect 12433 7712 12572 7714
rect 12433 7656 12438 7712
rect 12494 7656 12572 7712
rect 12433 7654 12572 7656
rect 12433 7651 12499 7654
rect 12566 7652 12572 7654
rect 12636 7652 12642 7716
rect 2646 7648 3042 7649
rect 2646 7584 2652 7648
rect 2716 7584 2732 7648
rect 2796 7584 2812 7648
rect 2876 7584 2892 7648
rect 2956 7584 2972 7648
rect 3036 7584 3042 7648
rect 2646 7583 3042 7584
rect 8646 7648 9042 7649
rect 8646 7584 8652 7648
rect 8716 7584 8732 7648
rect 8796 7584 8812 7648
rect 8876 7584 8892 7648
rect 8956 7584 8972 7648
rect 9036 7584 9042 7648
rect 8646 7583 9042 7584
rect 14646 7648 15042 7649
rect 14646 7584 14652 7648
rect 14716 7584 14732 7648
rect 14796 7584 14812 7648
rect 14876 7584 14892 7648
rect 14956 7584 14972 7648
rect 15036 7584 15042 7648
rect 14646 7583 15042 7584
rect 1906 7104 2302 7105
rect 1906 7040 1912 7104
rect 1976 7040 1992 7104
rect 2056 7040 2072 7104
rect 2136 7040 2152 7104
rect 2216 7040 2232 7104
rect 2296 7040 2302 7104
rect 1906 7039 2302 7040
rect 7906 7104 8302 7105
rect 7906 7040 7912 7104
rect 7976 7040 7992 7104
rect 8056 7040 8072 7104
rect 8136 7040 8152 7104
rect 8216 7040 8232 7104
rect 8296 7040 8302 7104
rect 7906 7039 8302 7040
rect 13906 7104 14302 7105
rect 13906 7040 13912 7104
rect 13976 7040 13992 7104
rect 14056 7040 14072 7104
rect 14136 7040 14152 7104
rect 14216 7040 14232 7104
rect 14296 7040 14302 7104
rect 13906 7039 14302 7040
rect 7833 6898 7899 6901
rect 14365 6898 14431 6901
rect 7833 6896 14431 6898
rect 7833 6840 7838 6896
rect 7894 6840 14370 6896
rect 14426 6840 14431 6896
rect 7833 6838 14431 6840
rect 7833 6835 7899 6838
rect 14365 6835 14431 6838
rect 7557 6762 7623 6765
rect 9397 6762 9463 6765
rect 7557 6760 9463 6762
rect 7557 6704 7562 6760
rect 7618 6704 9402 6760
rect 9458 6704 9463 6760
rect 7557 6702 9463 6704
rect 7557 6699 7623 6702
rect 9397 6699 9463 6702
rect 13445 6762 13511 6765
rect 13997 6762 14063 6765
rect 15561 6762 15627 6765
rect 13445 6760 15627 6762
rect 13445 6704 13450 6760
rect 13506 6704 14002 6760
rect 14058 6704 15566 6760
rect 15622 6704 15627 6760
rect 13445 6702 15627 6704
rect 13445 6699 13511 6702
rect 13997 6699 14063 6702
rect 15561 6699 15627 6702
rect 0 6626 800 6656
rect 1301 6626 1367 6629
rect 0 6624 1367 6626
rect 0 6568 1306 6624
rect 1362 6568 1367 6624
rect 0 6566 1367 6568
rect 0 6536 800 6566
rect 1301 6563 1367 6566
rect 2646 6560 3042 6561
rect 2646 6496 2652 6560
rect 2716 6496 2732 6560
rect 2796 6496 2812 6560
rect 2876 6496 2892 6560
rect 2956 6496 2972 6560
rect 3036 6496 3042 6560
rect 2646 6495 3042 6496
rect 8646 6560 9042 6561
rect 8646 6496 8652 6560
rect 8716 6496 8732 6560
rect 8796 6496 8812 6560
rect 8876 6496 8892 6560
rect 8956 6496 8972 6560
rect 9036 6496 9042 6560
rect 8646 6495 9042 6496
rect 14646 6560 15042 6561
rect 14646 6496 14652 6560
rect 14716 6496 14732 6560
rect 14796 6496 14812 6560
rect 14876 6496 14892 6560
rect 14956 6496 14972 6560
rect 15036 6496 15042 6560
rect 14646 6495 15042 6496
rect 14457 6492 14523 6493
rect 14406 6490 14412 6492
rect 14366 6430 14412 6490
rect 14476 6488 14523 6492
rect 14518 6432 14523 6488
rect 14406 6428 14412 6430
rect 14476 6428 14523 6432
rect 14457 6427 14523 6428
rect 6729 6354 6795 6357
rect 16481 6354 16547 6357
rect 6729 6352 16547 6354
rect 6729 6296 6734 6352
rect 6790 6296 16486 6352
rect 16542 6296 16547 6352
rect 6729 6294 16547 6296
rect 6729 6291 6795 6294
rect 16481 6291 16547 6294
rect 10685 6218 10751 6221
rect 16665 6218 16731 6221
rect 10685 6216 16731 6218
rect 10685 6160 10690 6216
rect 10746 6160 16670 6216
rect 16726 6160 16731 6216
rect 10685 6158 16731 6160
rect 10685 6155 10751 6158
rect 16665 6155 16731 6158
rect 1906 6016 2302 6017
rect 1906 5952 1912 6016
rect 1976 5952 1992 6016
rect 2056 5952 2072 6016
rect 2136 5952 2152 6016
rect 2216 5952 2232 6016
rect 2296 5952 2302 6016
rect 1906 5951 2302 5952
rect 7906 6016 8302 6017
rect 7906 5952 7912 6016
rect 7976 5952 7992 6016
rect 8056 5952 8072 6016
rect 8136 5952 8152 6016
rect 8216 5952 8232 6016
rect 8296 5952 8302 6016
rect 7906 5951 8302 5952
rect 13906 6016 14302 6017
rect 13906 5952 13912 6016
rect 13976 5952 13992 6016
rect 14056 5952 14072 6016
rect 14136 5952 14152 6016
rect 14216 5952 14232 6016
rect 14296 5952 14302 6016
rect 13906 5951 14302 5952
rect 0 5538 800 5568
rect 1393 5538 1459 5541
rect 0 5536 1459 5538
rect 0 5480 1398 5536
rect 1454 5480 1459 5536
rect 0 5478 1459 5480
rect 0 5448 800 5478
rect 1393 5475 1459 5478
rect 2646 5472 3042 5473
rect 2646 5408 2652 5472
rect 2716 5408 2732 5472
rect 2796 5408 2812 5472
rect 2876 5408 2892 5472
rect 2956 5408 2972 5472
rect 3036 5408 3042 5472
rect 2646 5407 3042 5408
rect 8646 5472 9042 5473
rect 8646 5408 8652 5472
rect 8716 5408 8732 5472
rect 8796 5408 8812 5472
rect 8876 5408 8892 5472
rect 8956 5408 8972 5472
rect 9036 5408 9042 5472
rect 8646 5407 9042 5408
rect 14646 5472 15042 5473
rect 14646 5408 14652 5472
rect 14716 5408 14732 5472
rect 14796 5408 14812 5472
rect 14876 5408 14892 5472
rect 14956 5408 14972 5472
rect 15036 5408 15042 5472
rect 14646 5407 15042 5408
rect 1906 4928 2302 4929
rect 1906 4864 1912 4928
rect 1976 4864 1992 4928
rect 2056 4864 2072 4928
rect 2136 4864 2152 4928
rect 2216 4864 2232 4928
rect 2296 4864 2302 4928
rect 1906 4863 2302 4864
rect 7906 4928 8302 4929
rect 7906 4864 7912 4928
rect 7976 4864 7992 4928
rect 8056 4864 8072 4928
rect 8136 4864 8152 4928
rect 8216 4864 8232 4928
rect 8296 4864 8302 4928
rect 7906 4863 8302 4864
rect 13906 4928 14302 4929
rect 13906 4864 13912 4928
rect 13976 4864 13992 4928
rect 14056 4864 14072 4928
rect 14136 4864 14152 4928
rect 14216 4864 14232 4928
rect 14296 4864 14302 4928
rect 13906 4863 14302 4864
rect 841 4586 907 4589
rect 798 4584 907 4586
rect 798 4528 846 4584
rect 902 4528 907 4584
rect 798 4523 907 4528
rect 798 4480 858 4523
rect 0 4390 858 4480
rect 0 4360 800 4390
rect 2646 4384 3042 4385
rect 2646 4320 2652 4384
rect 2716 4320 2732 4384
rect 2796 4320 2812 4384
rect 2876 4320 2892 4384
rect 2956 4320 2972 4384
rect 3036 4320 3042 4384
rect 2646 4319 3042 4320
rect 8646 4384 9042 4385
rect 8646 4320 8652 4384
rect 8716 4320 8732 4384
rect 8796 4320 8812 4384
rect 8876 4320 8892 4384
rect 8956 4320 8972 4384
rect 9036 4320 9042 4384
rect 8646 4319 9042 4320
rect 14646 4384 15042 4385
rect 14646 4320 14652 4384
rect 14716 4320 14732 4384
rect 14796 4320 14812 4384
rect 14876 4320 14892 4384
rect 14956 4320 14972 4384
rect 15036 4320 15042 4384
rect 14646 4319 15042 4320
rect 9765 4042 9831 4045
rect 11329 4042 11395 4045
rect 9765 4040 11395 4042
rect 9765 3984 9770 4040
rect 9826 3984 11334 4040
rect 11390 3984 11395 4040
rect 9765 3982 11395 3984
rect 9765 3979 9831 3982
rect 11329 3979 11395 3982
rect 1906 3840 2302 3841
rect 1906 3776 1912 3840
rect 1976 3776 1992 3840
rect 2056 3776 2072 3840
rect 2136 3776 2152 3840
rect 2216 3776 2232 3840
rect 2296 3776 2302 3840
rect 1906 3775 2302 3776
rect 7906 3840 8302 3841
rect 7906 3776 7912 3840
rect 7976 3776 7992 3840
rect 8056 3776 8072 3840
rect 8136 3776 8152 3840
rect 8216 3776 8232 3840
rect 8296 3776 8302 3840
rect 7906 3775 8302 3776
rect 13906 3840 14302 3841
rect 13906 3776 13912 3840
rect 13976 3776 13992 3840
rect 14056 3776 14072 3840
rect 14136 3776 14152 3840
rect 14216 3776 14232 3840
rect 14296 3776 14302 3840
rect 13906 3775 14302 3776
rect 841 3498 907 3501
rect 798 3496 907 3498
rect 798 3440 846 3496
rect 902 3440 907 3496
rect 798 3435 907 3440
rect 11605 3498 11671 3501
rect 15745 3498 15811 3501
rect 11605 3496 15811 3498
rect 11605 3440 11610 3496
rect 11666 3440 15750 3496
rect 15806 3440 15811 3496
rect 11605 3438 15811 3440
rect 11605 3435 11671 3438
rect 15745 3435 15811 3438
rect 798 3392 858 3435
rect 0 3302 858 3392
rect 0 3272 800 3302
rect 2646 3296 3042 3297
rect 2646 3232 2652 3296
rect 2716 3232 2732 3296
rect 2796 3232 2812 3296
rect 2876 3232 2892 3296
rect 2956 3232 2972 3296
rect 3036 3232 3042 3296
rect 2646 3231 3042 3232
rect 8646 3296 9042 3297
rect 8646 3232 8652 3296
rect 8716 3232 8732 3296
rect 8796 3232 8812 3296
rect 8876 3232 8892 3296
rect 8956 3232 8972 3296
rect 9036 3232 9042 3296
rect 8646 3231 9042 3232
rect 14646 3296 15042 3297
rect 14646 3232 14652 3296
rect 14716 3232 14732 3296
rect 14796 3232 14812 3296
rect 14876 3232 14892 3296
rect 14956 3232 14972 3296
rect 15036 3232 15042 3296
rect 14646 3231 15042 3232
rect 1906 2752 2302 2753
rect 1906 2688 1912 2752
rect 1976 2688 1992 2752
rect 2056 2688 2072 2752
rect 2136 2688 2152 2752
rect 2216 2688 2232 2752
rect 2296 2688 2302 2752
rect 1906 2687 2302 2688
rect 7906 2752 8302 2753
rect 7906 2688 7912 2752
rect 7976 2688 7992 2752
rect 8056 2688 8072 2752
rect 8136 2688 8152 2752
rect 8216 2688 8232 2752
rect 8296 2688 8302 2752
rect 7906 2687 8302 2688
rect 13906 2752 14302 2753
rect 13906 2688 13912 2752
rect 13976 2688 13992 2752
rect 14056 2688 14072 2752
rect 14136 2688 14152 2752
rect 14216 2688 14232 2752
rect 14296 2688 14302 2752
rect 13906 2687 14302 2688
rect 0 2274 800 2304
rect 1393 2274 1459 2277
rect 0 2272 1459 2274
rect 0 2216 1398 2272
rect 1454 2216 1459 2272
rect 0 2214 1459 2216
rect 0 2184 800 2214
rect 1393 2211 1459 2214
rect 2646 2208 3042 2209
rect 2646 2144 2652 2208
rect 2716 2144 2732 2208
rect 2796 2144 2812 2208
rect 2876 2144 2892 2208
rect 2956 2144 2972 2208
rect 3036 2144 3042 2208
rect 2646 2143 3042 2144
rect 8646 2208 9042 2209
rect 8646 2144 8652 2208
rect 8716 2144 8732 2208
rect 8796 2144 8812 2208
rect 8876 2144 8892 2208
rect 8956 2144 8972 2208
rect 9036 2144 9042 2208
rect 8646 2143 9042 2144
rect 14646 2208 15042 2209
rect 14646 2144 14652 2208
rect 14716 2144 14732 2208
rect 14796 2144 14812 2208
rect 14876 2144 14892 2208
rect 14956 2144 14972 2208
rect 15036 2144 15042 2208
rect 14646 2143 15042 2144
<< via3 >>
rect 2652 18524 2716 18528
rect 2652 18468 2656 18524
rect 2656 18468 2712 18524
rect 2712 18468 2716 18524
rect 2652 18464 2716 18468
rect 2732 18524 2796 18528
rect 2732 18468 2736 18524
rect 2736 18468 2792 18524
rect 2792 18468 2796 18524
rect 2732 18464 2796 18468
rect 2812 18524 2876 18528
rect 2812 18468 2816 18524
rect 2816 18468 2872 18524
rect 2872 18468 2876 18524
rect 2812 18464 2876 18468
rect 2892 18524 2956 18528
rect 2892 18468 2896 18524
rect 2896 18468 2952 18524
rect 2952 18468 2956 18524
rect 2892 18464 2956 18468
rect 2972 18524 3036 18528
rect 2972 18468 2976 18524
rect 2976 18468 3032 18524
rect 3032 18468 3036 18524
rect 2972 18464 3036 18468
rect 8652 18524 8716 18528
rect 8652 18468 8656 18524
rect 8656 18468 8712 18524
rect 8712 18468 8716 18524
rect 8652 18464 8716 18468
rect 8732 18524 8796 18528
rect 8732 18468 8736 18524
rect 8736 18468 8792 18524
rect 8792 18468 8796 18524
rect 8732 18464 8796 18468
rect 8812 18524 8876 18528
rect 8812 18468 8816 18524
rect 8816 18468 8872 18524
rect 8872 18468 8876 18524
rect 8812 18464 8876 18468
rect 8892 18524 8956 18528
rect 8892 18468 8896 18524
rect 8896 18468 8952 18524
rect 8952 18468 8956 18524
rect 8892 18464 8956 18468
rect 8972 18524 9036 18528
rect 8972 18468 8976 18524
rect 8976 18468 9032 18524
rect 9032 18468 9036 18524
rect 8972 18464 9036 18468
rect 14652 18524 14716 18528
rect 14652 18468 14656 18524
rect 14656 18468 14712 18524
rect 14712 18468 14716 18524
rect 14652 18464 14716 18468
rect 14732 18524 14796 18528
rect 14732 18468 14736 18524
rect 14736 18468 14792 18524
rect 14792 18468 14796 18524
rect 14732 18464 14796 18468
rect 14812 18524 14876 18528
rect 14812 18468 14816 18524
rect 14816 18468 14872 18524
rect 14872 18468 14876 18524
rect 14812 18464 14876 18468
rect 14892 18524 14956 18528
rect 14892 18468 14896 18524
rect 14896 18468 14952 18524
rect 14952 18468 14956 18524
rect 14892 18464 14956 18468
rect 14972 18524 15036 18528
rect 14972 18468 14976 18524
rect 14976 18468 15032 18524
rect 15032 18468 15036 18524
rect 14972 18464 15036 18468
rect 12572 17988 12636 18052
rect 1912 17980 1976 17984
rect 1912 17924 1916 17980
rect 1916 17924 1972 17980
rect 1972 17924 1976 17980
rect 1912 17920 1976 17924
rect 1992 17980 2056 17984
rect 1992 17924 1996 17980
rect 1996 17924 2052 17980
rect 2052 17924 2056 17980
rect 1992 17920 2056 17924
rect 2072 17980 2136 17984
rect 2072 17924 2076 17980
rect 2076 17924 2132 17980
rect 2132 17924 2136 17980
rect 2072 17920 2136 17924
rect 2152 17980 2216 17984
rect 2152 17924 2156 17980
rect 2156 17924 2212 17980
rect 2212 17924 2216 17980
rect 2152 17920 2216 17924
rect 2232 17980 2296 17984
rect 2232 17924 2236 17980
rect 2236 17924 2292 17980
rect 2292 17924 2296 17980
rect 2232 17920 2296 17924
rect 7912 17980 7976 17984
rect 7912 17924 7916 17980
rect 7916 17924 7972 17980
rect 7972 17924 7976 17980
rect 7912 17920 7976 17924
rect 7992 17980 8056 17984
rect 7992 17924 7996 17980
rect 7996 17924 8052 17980
rect 8052 17924 8056 17980
rect 7992 17920 8056 17924
rect 8072 17980 8136 17984
rect 8072 17924 8076 17980
rect 8076 17924 8132 17980
rect 8132 17924 8136 17980
rect 8072 17920 8136 17924
rect 8152 17980 8216 17984
rect 8152 17924 8156 17980
rect 8156 17924 8212 17980
rect 8212 17924 8216 17980
rect 8152 17920 8216 17924
rect 8232 17980 8296 17984
rect 8232 17924 8236 17980
rect 8236 17924 8292 17980
rect 8292 17924 8296 17980
rect 8232 17920 8296 17924
rect 13912 17980 13976 17984
rect 13912 17924 13916 17980
rect 13916 17924 13972 17980
rect 13972 17924 13976 17980
rect 13912 17920 13976 17924
rect 13992 17980 14056 17984
rect 13992 17924 13996 17980
rect 13996 17924 14052 17980
rect 14052 17924 14056 17980
rect 13992 17920 14056 17924
rect 14072 17980 14136 17984
rect 14072 17924 14076 17980
rect 14076 17924 14132 17980
rect 14132 17924 14136 17980
rect 14072 17920 14136 17924
rect 14152 17980 14216 17984
rect 14152 17924 14156 17980
rect 14156 17924 14212 17980
rect 14212 17924 14216 17980
rect 14152 17920 14216 17924
rect 14232 17980 14296 17984
rect 14232 17924 14236 17980
rect 14236 17924 14292 17980
rect 14292 17924 14296 17980
rect 14232 17920 14296 17924
rect 2652 17436 2716 17440
rect 2652 17380 2656 17436
rect 2656 17380 2712 17436
rect 2712 17380 2716 17436
rect 2652 17376 2716 17380
rect 2732 17436 2796 17440
rect 2732 17380 2736 17436
rect 2736 17380 2792 17436
rect 2792 17380 2796 17436
rect 2732 17376 2796 17380
rect 2812 17436 2876 17440
rect 2812 17380 2816 17436
rect 2816 17380 2872 17436
rect 2872 17380 2876 17436
rect 2812 17376 2876 17380
rect 2892 17436 2956 17440
rect 2892 17380 2896 17436
rect 2896 17380 2952 17436
rect 2952 17380 2956 17436
rect 2892 17376 2956 17380
rect 2972 17436 3036 17440
rect 2972 17380 2976 17436
rect 2976 17380 3032 17436
rect 3032 17380 3036 17436
rect 2972 17376 3036 17380
rect 8652 17436 8716 17440
rect 8652 17380 8656 17436
rect 8656 17380 8712 17436
rect 8712 17380 8716 17436
rect 8652 17376 8716 17380
rect 8732 17436 8796 17440
rect 8732 17380 8736 17436
rect 8736 17380 8792 17436
rect 8792 17380 8796 17436
rect 8732 17376 8796 17380
rect 8812 17436 8876 17440
rect 8812 17380 8816 17436
rect 8816 17380 8872 17436
rect 8872 17380 8876 17436
rect 8812 17376 8876 17380
rect 8892 17436 8956 17440
rect 8892 17380 8896 17436
rect 8896 17380 8952 17436
rect 8952 17380 8956 17436
rect 8892 17376 8956 17380
rect 8972 17436 9036 17440
rect 8972 17380 8976 17436
rect 8976 17380 9032 17436
rect 9032 17380 9036 17436
rect 8972 17376 9036 17380
rect 14652 17436 14716 17440
rect 14652 17380 14656 17436
rect 14656 17380 14712 17436
rect 14712 17380 14716 17436
rect 14652 17376 14716 17380
rect 14732 17436 14796 17440
rect 14732 17380 14736 17436
rect 14736 17380 14792 17436
rect 14792 17380 14796 17436
rect 14732 17376 14796 17380
rect 14812 17436 14876 17440
rect 14812 17380 14816 17436
rect 14816 17380 14872 17436
rect 14872 17380 14876 17436
rect 14812 17376 14876 17380
rect 14892 17436 14956 17440
rect 14892 17380 14896 17436
rect 14896 17380 14952 17436
rect 14952 17380 14956 17436
rect 14892 17376 14956 17380
rect 14972 17436 15036 17440
rect 14972 17380 14976 17436
rect 14976 17380 15032 17436
rect 15032 17380 15036 17436
rect 14972 17376 15036 17380
rect 1912 16892 1976 16896
rect 1912 16836 1916 16892
rect 1916 16836 1972 16892
rect 1972 16836 1976 16892
rect 1912 16832 1976 16836
rect 1992 16892 2056 16896
rect 1992 16836 1996 16892
rect 1996 16836 2052 16892
rect 2052 16836 2056 16892
rect 1992 16832 2056 16836
rect 2072 16892 2136 16896
rect 2072 16836 2076 16892
rect 2076 16836 2132 16892
rect 2132 16836 2136 16892
rect 2072 16832 2136 16836
rect 2152 16892 2216 16896
rect 2152 16836 2156 16892
rect 2156 16836 2212 16892
rect 2212 16836 2216 16892
rect 2152 16832 2216 16836
rect 2232 16892 2296 16896
rect 2232 16836 2236 16892
rect 2236 16836 2292 16892
rect 2292 16836 2296 16892
rect 2232 16832 2296 16836
rect 7912 16892 7976 16896
rect 7912 16836 7916 16892
rect 7916 16836 7972 16892
rect 7972 16836 7976 16892
rect 7912 16832 7976 16836
rect 7992 16892 8056 16896
rect 7992 16836 7996 16892
rect 7996 16836 8052 16892
rect 8052 16836 8056 16892
rect 7992 16832 8056 16836
rect 8072 16892 8136 16896
rect 8072 16836 8076 16892
rect 8076 16836 8132 16892
rect 8132 16836 8136 16892
rect 8072 16832 8136 16836
rect 8152 16892 8216 16896
rect 8152 16836 8156 16892
rect 8156 16836 8212 16892
rect 8212 16836 8216 16892
rect 8152 16832 8216 16836
rect 8232 16892 8296 16896
rect 8232 16836 8236 16892
rect 8236 16836 8292 16892
rect 8292 16836 8296 16892
rect 8232 16832 8296 16836
rect 13912 16892 13976 16896
rect 13912 16836 13916 16892
rect 13916 16836 13972 16892
rect 13972 16836 13976 16892
rect 13912 16832 13976 16836
rect 13992 16892 14056 16896
rect 13992 16836 13996 16892
rect 13996 16836 14052 16892
rect 14052 16836 14056 16892
rect 13992 16832 14056 16836
rect 14072 16892 14136 16896
rect 14072 16836 14076 16892
rect 14076 16836 14132 16892
rect 14132 16836 14136 16892
rect 14072 16832 14136 16836
rect 14152 16892 14216 16896
rect 14152 16836 14156 16892
rect 14156 16836 14212 16892
rect 14212 16836 14216 16892
rect 14152 16832 14216 16836
rect 14232 16892 14296 16896
rect 14232 16836 14236 16892
rect 14236 16836 14292 16892
rect 14292 16836 14296 16892
rect 14232 16832 14296 16836
rect 2652 16348 2716 16352
rect 2652 16292 2656 16348
rect 2656 16292 2712 16348
rect 2712 16292 2716 16348
rect 2652 16288 2716 16292
rect 2732 16348 2796 16352
rect 2732 16292 2736 16348
rect 2736 16292 2792 16348
rect 2792 16292 2796 16348
rect 2732 16288 2796 16292
rect 2812 16348 2876 16352
rect 2812 16292 2816 16348
rect 2816 16292 2872 16348
rect 2872 16292 2876 16348
rect 2812 16288 2876 16292
rect 2892 16348 2956 16352
rect 2892 16292 2896 16348
rect 2896 16292 2952 16348
rect 2952 16292 2956 16348
rect 2892 16288 2956 16292
rect 2972 16348 3036 16352
rect 2972 16292 2976 16348
rect 2976 16292 3032 16348
rect 3032 16292 3036 16348
rect 2972 16288 3036 16292
rect 8652 16348 8716 16352
rect 8652 16292 8656 16348
rect 8656 16292 8712 16348
rect 8712 16292 8716 16348
rect 8652 16288 8716 16292
rect 8732 16348 8796 16352
rect 8732 16292 8736 16348
rect 8736 16292 8792 16348
rect 8792 16292 8796 16348
rect 8732 16288 8796 16292
rect 8812 16348 8876 16352
rect 8812 16292 8816 16348
rect 8816 16292 8872 16348
rect 8872 16292 8876 16348
rect 8812 16288 8876 16292
rect 8892 16348 8956 16352
rect 8892 16292 8896 16348
rect 8896 16292 8952 16348
rect 8952 16292 8956 16348
rect 8892 16288 8956 16292
rect 8972 16348 9036 16352
rect 8972 16292 8976 16348
rect 8976 16292 9032 16348
rect 9032 16292 9036 16348
rect 8972 16288 9036 16292
rect 14652 16348 14716 16352
rect 14652 16292 14656 16348
rect 14656 16292 14712 16348
rect 14712 16292 14716 16348
rect 14652 16288 14716 16292
rect 14732 16348 14796 16352
rect 14732 16292 14736 16348
rect 14736 16292 14792 16348
rect 14792 16292 14796 16348
rect 14732 16288 14796 16292
rect 14812 16348 14876 16352
rect 14812 16292 14816 16348
rect 14816 16292 14872 16348
rect 14872 16292 14876 16348
rect 14812 16288 14876 16292
rect 14892 16348 14956 16352
rect 14892 16292 14896 16348
rect 14896 16292 14952 16348
rect 14952 16292 14956 16348
rect 14892 16288 14956 16292
rect 14972 16348 15036 16352
rect 14972 16292 14976 16348
rect 14976 16292 15032 16348
rect 15032 16292 15036 16348
rect 14972 16288 15036 16292
rect 1912 15804 1976 15808
rect 1912 15748 1916 15804
rect 1916 15748 1972 15804
rect 1972 15748 1976 15804
rect 1912 15744 1976 15748
rect 1992 15804 2056 15808
rect 1992 15748 1996 15804
rect 1996 15748 2052 15804
rect 2052 15748 2056 15804
rect 1992 15744 2056 15748
rect 2072 15804 2136 15808
rect 2072 15748 2076 15804
rect 2076 15748 2132 15804
rect 2132 15748 2136 15804
rect 2072 15744 2136 15748
rect 2152 15804 2216 15808
rect 2152 15748 2156 15804
rect 2156 15748 2212 15804
rect 2212 15748 2216 15804
rect 2152 15744 2216 15748
rect 2232 15804 2296 15808
rect 2232 15748 2236 15804
rect 2236 15748 2292 15804
rect 2292 15748 2296 15804
rect 2232 15744 2296 15748
rect 7912 15804 7976 15808
rect 7912 15748 7916 15804
rect 7916 15748 7972 15804
rect 7972 15748 7976 15804
rect 7912 15744 7976 15748
rect 7992 15804 8056 15808
rect 7992 15748 7996 15804
rect 7996 15748 8052 15804
rect 8052 15748 8056 15804
rect 7992 15744 8056 15748
rect 8072 15804 8136 15808
rect 8072 15748 8076 15804
rect 8076 15748 8132 15804
rect 8132 15748 8136 15804
rect 8072 15744 8136 15748
rect 8152 15804 8216 15808
rect 8152 15748 8156 15804
rect 8156 15748 8212 15804
rect 8212 15748 8216 15804
rect 8152 15744 8216 15748
rect 8232 15804 8296 15808
rect 8232 15748 8236 15804
rect 8236 15748 8292 15804
rect 8292 15748 8296 15804
rect 8232 15744 8296 15748
rect 13912 15804 13976 15808
rect 13912 15748 13916 15804
rect 13916 15748 13972 15804
rect 13972 15748 13976 15804
rect 13912 15744 13976 15748
rect 13992 15804 14056 15808
rect 13992 15748 13996 15804
rect 13996 15748 14052 15804
rect 14052 15748 14056 15804
rect 13992 15744 14056 15748
rect 14072 15804 14136 15808
rect 14072 15748 14076 15804
rect 14076 15748 14132 15804
rect 14132 15748 14136 15804
rect 14072 15744 14136 15748
rect 14152 15804 14216 15808
rect 14152 15748 14156 15804
rect 14156 15748 14212 15804
rect 14212 15748 14216 15804
rect 14152 15744 14216 15748
rect 14232 15804 14296 15808
rect 14232 15748 14236 15804
rect 14236 15748 14292 15804
rect 14292 15748 14296 15804
rect 14232 15744 14296 15748
rect 2652 15260 2716 15264
rect 2652 15204 2656 15260
rect 2656 15204 2712 15260
rect 2712 15204 2716 15260
rect 2652 15200 2716 15204
rect 2732 15260 2796 15264
rect 2732 15204 2736 15260
rect 2736 15204 2792 15260
rect 2792 15204 2796 15260
rect 2732 15200 2796 15204
rect 2812 15260 2876 15264
rect 2812 15204 2816 15260
rect 2816 15204 2872 15260
rect 2872 15204 2876 15260
rect 2812 15200 2876 15204
rect 2892 15260 2956 15264
rect 2892 15204 2896 15260
rect 2896 15204 2952 15260
rect 2952 15204 2956 15260
rect 2892 15200 2956 15204
rect 2972 15260 3036 15264
rect 2972 15204 2976 15260
rect 2976 15204 3032 15260
rect 3032 15204 3036 15260
rect 2972 15200 3036 15204
rect 8652 15260 8716 15264
rect 8652 15204 8656 15260
rect 8656 15204 8712 15260
rect 8712 15204 8716 15260
rect 8652 15200 8716 15204
rect 8732 15260 8796 15264
rect 8732 15204 8736 15260
rect 8736 15204 8792 15260
rect 8792 15204 8796 15260
rect 8732 15200 8796 15204
rect 8812 15260 8876 15264
rect 8812 15204 8816 15260
rect 8816 15204 8872 15260
rect 8872 15204 8876 15260
rect 8812 15200 8876 15204
rect 8892 15260 8956 15264
rect 8892 15204 8896 15260
rect 8896 15204 8952 15260
rect 8952 15204 8956 15260
rect 8892 15200 8956 15204
rect 8972 15260 9036 15264
rect 8972 15204 8976 15260
rect 8976 15204 9032 15260
rect 9032 15204 9036 15260
rect 8972 15200 9036 15204
rect 14652 15260 14716 15264
rect 14652 15204 14656 15260
rect 14656 15204 14712 15260
rect 14712 15204 14716 15260
rect 14652 15200 14716 15204
rect 14732 15260 14796 15264
rect 14732 15204 14736 15260
rect 14736 15204 14792 15260
rect 14792 15204 14796 15260
rect 14732 15200 14796 15204
rect 14812 15260 14876 15264
rect 14812 15204 14816 15260
rect 14816 15204 14872 15260
rect 14872 15204 14876 15260
rect 14812 15200 14876 15204
rect 14892 15260 14956 15264
rect 14892 15204 14896 15260
rect 14896 15204 14952 15260
rect 14952 15204 14956 15260
rect 14892 15200 14956 15204
rect 14972 15260 15036 15264
rect 14972 15204 14976 15260
rect 14976 15204 15032 15260
rect 15032 15204 15036 15260
rect 14972 15200 15036 15204
rect 1912 14716 1976 14720
rect 1912 14660 1916 14716
rect 1916 14660 1972 14716
rect 1972 14660 1976 14716
rect 1912 14656 1976 14660
rect 1992 14716 2056 14720
rect 1992 14660 1996 14716
rect 1996 14660 2052 14716
rect 2052 14660 2056 14716
rect 1992 14656 2056 14660
rect 2072 14716 2136 14720
rect 2072 14660 2076 14716
rect 2076 14660 2132 14716
rect 2132 14660 2136 14716
rect 2072 14656 2136 14660
rect 2152 14716 2216 14720
rect 2152 14660 2156 14716
rect 2156 14660 2212 14716
rect 2212 14660 2216 14716
rect 2152 14656 2216 14660
rect 2232 14716 2296 14720
rect 2232 14660 2236 14716
rect 2236 14660 2292 14716
rect 2292 14660 2296 14716
rect 2232 14656 2296 14660
rect 7912 14716 7976 14720
rect 7912 14660 7916 14716
rect 7916 14660 7972 14716
rect 7972 14660 7976 14716
rect 7912 14656 7976 14660
rect 7992 14716 8056 14720
rect 7992 14660 7996 14716
rect 7996 14660 8052 14716
rect 8052 14660 8056 14716
rect 7992 14656 8056 14660
rect 8072 14716 8136 14720
rect 8072 14660 8076 14716
rect 8076 14660 8132 14716
rect 8132 14660 8136 14716
rect 8072 14656 8136 14660
rect 8152 14716 8216 14720
rect 8152 14660 8156 14716
rect 8156 14660 8212 14716
rect 8212 14660 8216 14716
rect 8152 14656 8216 14660
rect 8232 14716 8296 14720
rect 8232 14660 8236 14716
rect 8236 14660 8292 14716
rect 8292 14660 8296 14716
rect 8232 14656 8296 14660
rect 13912 14716 13976 14720
rect 13912 14660 13916 14716
rect 13916 14660 13972 14716
rect 13972 14660 13976 14716
rect 13912 14656 13976 14660
rect 13992 14716 14056 14720
rect 13992 14660 13996 14716
rect 13996 14660 14052 14716
rect 14052 14660 14056 14716
rect 13992 14656 14056 14660
rect 14072 14716 14136 14720
rect 14072 14660 14076 14716
rect 14076 14660 14132 14716
rect 14132 14660 14136 14716
rect 14072 14656 14136 14660
rect 14152 14716 14216 14720
rect 14152 14660 14156 14716
rect 14156 14660 14212 14716
rect 14212 14660 14216 14716
rect 14152 14656 14216 14660
rect 14232 14716 14296 14720
rect 14232 14660 14236 14716
rect 14236 14660 14292 14716
rect 14292 14660 14296 14716
rect 14232 14656 14296 14660
rect 2652 14172 2716 14176
rect 2652 14116 2656 14172
rect 2656 14116 2712 14172
rect 2712 14116 2716 14172
rect 2652 14112 2716 14116
rect 2732 14172 2796 14176
rect 2732 14116 2736 14172
rect 2736 14116 2792 14172
rect 2792 14116 2796 14172
rect 2732 14112 2796 14116
rect 2812 14172 2876 14176
rect 2812 14116 2816 14172
rect 2816 14116 2872 14172
rect 2872 14116 2876 14172
rect 2812 14112 2876 14116
rect 2892 14172 2956 14176
rect 2892 14116 2896 14172
rect 2896 14116 2952 14172
rect 2952 14116 2956 14172
rect 2892 14112 2956 14116
rect 2972 14172 3036 14176
rect 2972 14116 2976 14172
rect 2976 14116 3032 14172
rect 3032 14116 3036 14172
rect 2972 14112 3036 14116
rect 8652 14172 8716 14176
rect 8652 14116 8656 14172
rect 8656 14116 8712 14172
rect 8712 14116 8716 14172
rect 8652 14112 8716 14116
rect 8732 14172 8796 14176
rect 8732 14116 8736 14172
rect 8736 14116 8792 14172
rect 8792 14116 8796 14172
rect 8732 14112 8796 14116
rect 8812 14172 8876 14176
rect 8812 14116 8816 14172
rect 8816 14116 8872 14172
rect 8872 14116 8876 14172
rect 8812 14112 8876 14116
rect 8892 14172 8956 14176
rect 8892 14116 8896 14172
rect 8896 14116 8952 14172
rect 8952 14116 8956 14172
rect 8892 14112 8956 14116
rect 8972 14172 9036 14176
rect 8972 14116 8976 14172
rect 8976 14116 9032 14172
rect 9032 14116 9036 14172
rect 8972 14112 9036 14116
rect 14652 14172 14716 14176
rect 14652 14116 14656 14172
rect 14656 14116 14712 14172
rect 14712 14116 14716 14172
rect 14652 14112 14716 14116
rect 14732 14172 14796 14176
rect 14732 14116 14736 14172
rect 14736 14116 14792 14172
rect 14792 14116 14796 14172
rect 14732 14112 14796 14116
rect 14812 14172 14876 14176
rect 14812 14116 14816 14172
rect 14816 14116 14872 14172
rect 14872 14116 14876 14172
rect 14812 14112 14876 14116
rect 14892 14172 14956 14176
rect 14892 14116 14896 14172
rect 14896 14116 14952 14172
rect 14952 14116 14956 14172
rect 14892 14112 14956 14116
rect 14972 14172 15036 14176
rect 14972 14116 14976 14172
rect 14976 14116 15032 14172
rect 15032 14116 15036 14172
rect 14972 14112 15036 14116
rect 1912 13628 1976 13632
rect 1912 13572 1916 13628
rect 1916 13572 1972 13628
rect 1972 13572 1976 13628
rect 1912 13568 1976 13572
rect 1992 13628 2056 13632
rect 1992 13572 1996 13628
rect 1996 13572 2052 13628
rect 2052 13572 2056 13628
rect 1992 13568 2056 13572
rect 2072 13628 2136 13632
rect 2072 13572 2076 13628
rect 2076 13572 2132 13628
rect 2132 13572 2136 13628
rect 2072 13568 2136 13572
rect 2152 13628 2216 13632
rect 2152 13572 2156 13628
rect 2156 13572 2212 13628
rect 2212 13572 2216 13628
rect 2152 13568 2216 13572
rect 2232 13628 2296 13632
rect 2232 13572 2236 13628
rect 2236 13572 2292 13628
rect 2292 13572 2296 13628
rect 2232 13568 2296 13572
rect 7912 13628 7976 13632
rect 7912 13572 7916 13628
rect 7916 13572 7972 13628
rect 7972 13572 7976 13628
rect 7912 13568 7976 13572
rect 7992 13628 8056 13632
rect 7992 13572 7996 13628
rect 7996 13572 8052 13628
rect 8052 13572 8056 13628
rect 7992 13568 8056 13572
rect 8072 13628 8136 13632
rect 8072 13572 8076 13628
rect 8076 13572 8132 13628
rect 8132 13572 8136 13628
rect 8072 13568 8136 13572
rect 8152 13628 8216 13632
rect 8152 13572 8156 13628
rect 8156 13572 8212 13628
rect 8212 13572 8216 13628
rect 8152 13568 8216 13572
rect 8232 13628 8296 13632
rect 8232 13572 8236 13628
rect 8236 13572 8292 13628
rect 8292 13572 8296 13628
rect 8232 13568 8296 13572
rect 13912 13628 13976 13632
rect 13912 13572 13916 13628
rect 13916 13572 13972 13628
rect 13972 13572 13976 13628
rect 13912 13568 13976 13572
rect 13992 13628 14056 13632
rect 13992 13572 13996 13628
rect 13996 13572 14052 13628
rect 14052 13572 14056 13628
rect 13992 13568 14056 13572
rect 14072 13628 14136 13632
rect 14072 13572 14076 13628
rect 14076 13572 14132 13628
rect 14132 13572 14136 13628
rect 14072 13568 14136 13572
rect 14152 13628 14216 13632
rect 14152 13572 14156 13628
rect 14156 13572 14212 13628
rect 14212 13572 14216 13628
rect 14152 13568 14216 13572
rect 14232 13628 14296 13632
rect 14232 13572 14236 13628
rect 14236 13572 14292 13628
rect 14292 13572 14296 13628
rect 14232 13568 14296 13572
rect 2652 13084 2716 13088
rect 2652 13028 2656 13084
rect 2656 13028 2712 13084
rect 2712 13028 2716 13084
rect 2652 13024 2716 13028
rect 2732 13084 2796 13088
rect 2732 13028 2736 13084
rect 2736 13028 2792 13084
rect 2792 13028 2796 13084
rect 2732 13024 2796 13028
rect 2812 13084 2876 13088
rect 2812 13028 2816 13084
rect 2816 13028 2872 13084
rect 2872 13028 2876 13084
rect 2812 13024 2876 13028
rect 2892 13084 2956 13088
rect 2892 13028 2896 13084
rect 2896 13028 2952 13084
rect 2952 13028 2956 13084
rect 2892 13024 2956 13028
rect 2972 13084 3036 13088
rect 2972 13028 2976 13084
rect 2976 13028 3032 13084
rect 3032 13028 3036 13084
rect 2972 13024 3036 13028
rect 8652 13084 8716 13088
rect 8652 13028 8656 13084
rect 8656 13028 8712 13084
rect 8712 13028 8716 13084
rect 8652 13024 8716 13028
rect 8732 13084 8796 13088
rect 8732 13028 8736 13084
rect 8736 13028 8792 13084
rect 8792 13028 8796 13084
rect 8732 13024 8796 13028
rect 8812 13084 8876 13088
rect 8812 13028 8816 13084
rect 8816 13028 8872 13084
rect 8872 13028 8876 13084
rect 8812 13024 8876 13028
rect 8892 13084 8956 13088
rect 8892 13028 8896 13084
rect 8896 13028 8952 13084
rect 8952 13028 8956 13084
rect 8892 13024 8956 13028
rect 8972 13084 9036 13088
rect 8972 13028 8976 13084
rect 8976 13028 9032 13084
rect 9032 13028 9036 13084
rect 8972 13024 9036 13028
rect 14652 13084 14716 13088
rect 14652 13028 14656 13084
rect 14656 13028 14712 13084
rect 14712 13028 14716 13084
rect 14652 13024 14716 13028
rect 14732 13084 14796 13088
rect 14732 13028 14736 13084
rect 14736 13028 14792 13084
rect 14792 13028 14796 13084
rect 14732 13024 14796 13028
rect 14812 13084 14876 13088
rect 14812 13028 14816 13084
rect 14816 13028 14872 13084
rect 14872 13028 14876 13084
rect 14812 13024 14876 13028
rect 14892 13084 14956 13088
rect 14892 13028 14896 13084
rect 14896 13028 14952 13084
rect 14952 13028 14956 13084
rect 14892 13024 14956 13028
rect 14972 13084 15036 13088
rect 14972 13028 14976 13084
rect 14976 13028 15032 13084
rect 15032 13028 15036 13084
rect 14972 13024 15036 13028
rect 1912 12540 1976 12544
rect 1912 12484 1916 12540
rect 1916 12484 1972 12540
rect 1972 12484 1976 12540
rect 1912 12480 1976 12484
rect 1992 12540 2056 12544
rect 1992 12484 1996 12540
rect 1996 12484 2052 12540
rect 2052 12484 2056 12540
rect 1992 12480 2056 12484
rect 2072 12540 2136 12544
rect 2072 12484 2076 12540
rect 2076 12484 2132 12540
rect 2132 12484 2136 12540
rect 2072 12480 2136 12484
rect 2152 12540 2216 12544
rect 2152 12484 2156 12540
rect 2156 12484 2212 12540
rect 2212 12484 2216 12540
rect 2152 12480 2216 12484
rect 2232 12540 2296 12544
rect 2232 12484 2236 12540
rect 2236 12484 2292 12540
rect 2292 12484 2296 12540
rect 2232 12480 2296 12484
rect 7912 12540 7976 12544
rect 7912 12484 7916 12540
rect 7916 12484 7972 12540
rect 7972 12484 7976 12540
rect 7912 12480 7976 12484
rect 7992 12540 8056 12544
rect 7992 12484 7996 12540
rect 7996 12484 8052 12540
rect 8052 12484 8056 12540
rect 7992 12480 8056 12484
rect 8072 12540 8136 12544
rect 8072 12484 8076 12540
rect 8076 12484 8132 12540
rect 8132 12484 8136 12540
rect 8072 12480 8136 12484
rect 8152 12540 8216 12544
rect 8152 12484 8156 12540
rect 8156 12484 8212 12540
rect 8212 12484 8216 12540
rect 8152 12480 8216 12484
rect 8232 12540 8296 12544
rect 8232 12484 8236 12540
rect 8236 12484 8292 12540
rect 8292 12484 8296 12540
rect 8232 12480 8296 12484
rect 13912 12540 13976 12544
rect 13912 12484 13916 12540
rect 13916 12484 13972 12540
rect 13972 12484 13976 12540
rect 13912 12480 13976 12484
rect 13992 12540 14056 12544
rect 13992 12484 13996 12540
rect 13996 12484 14052 12540
rect 14052 12484 14056 12540
rect 13992 12480 14056 12484
rect 14072 12540 14136 12544
rect 14072 12484 14076 12540
rect 14076 12484 14132 12540
rect 14132 12484 14136 12540
rect 14072 12480 14136 12484
rect 14152 12540 14216 12544
rect 14152 12484 14156 12540
rect 14156 12484 14212 12540
rect 14212 12484 14216 12540
rect 14152 12480 14216 12484
rect 14232 12540 14296 12544
rect 14232 12484 14236 12540
rect 14236 12484 14292 12540
rect 14292 12484 14296 12540
rect 14232 12480 14296 12484
rect 2652 11996 2716 12000
rect 2652 11940 2656 11996
rect 2656 11940 2712 11996
rect 2712 11940 2716 11996
rect 2652 11936 2716 11940
rect 2732 11996 2796 12000
rect 2732 11940 2736 11996
rect 2736 11940 2792 11996
rect 2792 11940 2796 11996
rect 2732 11936 2796 11940
rect 2812 11996 2876 12000
rect 2812 11940 2816 11996
rect 2816 11940 2872 11996
rect 2872 11940 2876 11996
rect 2812 11936 2876 11940
rect 2892 11996 2956 12000
rect 2892 11940 2896 11996
rect 2896 11940 2952 11996
rect 2952 11940 2956 11996
rect 2892 11936 2956 11940
rect 2972 11996 3036 12000
rect 2972 11940 2976 11996
rect 2976 11940 3032 11996
rect 3032 11940 3036 11996
rect 2972 11936 3036 11940
rect 8652 11996 8716 12000
rect 8652 11940 8656 11996
rect 8656 11940 8712 11996
rect 8712 11940 8716 11996
rect 8652 11936 8716 11940
rect 8732 11996 8796 12000
rect 8732 11940 8736 11996
rect 8736 11940 8792 11996
rect 8792 11940 8796 11996
rect 8732 11936 8796 11940
rect 8812 11996 8876 12000
rect 8812 11940 8816 11996
rect 8816 11940 8872 11996
rect 8872 11940 8876 11996
rect 8812 11936 8876 11940
rect 8892 11996 8956 12000
rect 8892 11940 8896 11996
rect 8896 11940 8952 11996
rect 8952 11940 8956 11996
rect 8892 11936 8956 11940
rect 8972 11996 9036 12000
rect 8972 11940 8976 11996
rect 8976 11940 9032 11996
rect 9032 11940 9036 11996
rect 8972 11936 9036 11940
rect 14652 11996 14716 12000
rect 14652 11940 14656 11996
rect 14656 11940 14712 11996
rect 14712 11940 14716 11996
rect 14652 11936 14716 11940
rect 14732 11996 14796 12000
rect 14732 11940 14736 11996
rect 14736 11940 14792 11996
rect 14792 11940 14796 11996
rect 14732 11936 14796 11940
rect 14812 11996 14876 12000
rect 14812 11940 14816 11996
rect 14816 11940 14872 11996
rect 14872 11940 14876 11996
rect 14812 11936 14876 11940
rect 14892 11996 14956 12000
rect 14892 11940 14896 11996
rect 14896 11940 14952 11996
rect 14952 11940 14956 11996
rect 14892 11936 14956 11940
rect 14972 11996 15036 12000
rect 14972 11940 14976 11996
rect 14976 11940 15032 11996
rect 15032 11940 15036 11996
rect 14972 11936 15036 11940
rect 1912 11452 1976 11456
rect 1912 11396 1916 11452
rect 1916 11396 1972 11452
rect 1972 11396 1976 11452
rect 1912 11392 1976 11396
rect 1992 11452 2056 11456
rect 1992 11396 1996 11452
rect 1996 11396 2052 11452
rect 2052 11396 2056 11452
rect 1992 11392 2056 11396
rect 2072 11452 2136 11456
rect 2072 11396 2076 11452
rect 2076 11396 2132 11452
rect 2132 11396 2136 11452
rect 2072 11392 2136 11396
rect 2152 11452 2216 11456
rect 2152 11396 2156 11452
rect 2156 11396 2212 11452
rect 2212 11396 2216 11452
rect 2152 11392 2216 11396
rect 2232 11452 2296 11456
rect 2232 11396 2236 11452
rect 2236 11396 2292 11452
rect 2292 11396 2296 11452
rect 2232 11392 2296 11396
rect 7912 11452 7976 11456
rect 7912 11396 7916 11452
rect 7916 11396 7972 11452
rect 7972 11396 7976 11452
rect 7912 11392 7976 11396
rect 7992 11452 8056 11456
rect 7992 11396 7996 11452
rect 7996 11396 8052 11452
rect 8052 11396 8056 11452
rect 7992 11392 8056 11396
rect 8072 11452 8136 11456
rect 8072 11396 8076 11452
rect 8076 11396 8132 11452
rect 8132 11396 8136 11452
rect 8072 11392 8136 11396
rect 8152 11452 8216 11456
rect 8152 11396 8156 11452
rect 8156 11396 8212 11452
rect 8212 11396 8216 11452
rect 8152 11392 8216 11396
rect 8232 11452 8296 11456
rect 8232 11396 8236 11452
rect 8236 11396 8292 11452
rect 8292 11396 8296 11452
rect 8232 11392 8296 11396
rect 13912 11452 13976 11456
rect 13912 11396 13916 11452
rect 13916 11396 13972 11452
rect 13972 11396 13976 11452
rect 13912 11392 13976 11396
rect 13992 11452 14056 11456
rect 13992 11396 13996 11452
rect 13996 11396 14052 11452
rect 14052 11396 14056 11452
rect 13992 11392 14056 11396
rect 14072 11452 14136 11456
rect 14072 11396 14076 11452
rect 14076 11396 14132 11452
rect 14132 11396 14136 11452
rect 14072 11392 14136 11396
rect 14152 11452 14216 11456
rect 14152 11396 14156 11452
rect 14156 11396 14212 11452
rect 14212 11396 14216 11452
rect 14152 11392 14216 11396
rect 14232 11452 14296 11456
rect 14232 11396 14236 11452
rect 14236 11396 14292 11452
rect 14292 11396 14296 11452
rect 14232 11392 14296 11396
rect 2652 10908 2716 10912
rect 2652 10852 2656 10908
rect 2656 10852 2712 10908
rect 2712 10852 2716 10908
rect 2652 10848 2716 10852
rect 2732 10908 2796 10912
rect 2732 10852 2736 10908
rect 2736 10852 2792 10908
rect 2792 10852 2796 10908
rect 2732 10848 2796 10852
rect 2812 10908 2876 10912
rect 2812 10852 2816 10908
rect 2816 10852 2872 10908
rect 2872 10852 2876 10908
rect 2812 10848 2876 10852
rect 2892 10908 2956 10912
rect 2892 10852 2896 10908
rect 2896 10852 2952 10908
rect 2952 10852 2956 10908
rect 2892 10848 2956 10852
rect 2972 10908 3036 10912
rect 2972 10852 2976 10908
rect 2976 10852 3032 10908
rect 3032 10852 3036 10908
rect 2972 10848 3036 10852
rect 8652 10908 8716 10912
rect 8652 10852 8656 10908
rect 8656 10852 8712 10908
rect 8712 10852 8716 10908
rect 8652 10848 8716 10852
rect 8732 10908 8796 10912
rect 8732 10852 8736 10908
rect 8736 10852 8792 10908
rect 8792 10852 8796 10908
rect 8732 10848 8796 10852
rect 8812 10908 8876 10912
rect 8812 10852 8816 10908
rect 8816 10852 8872 10908
rect 8872 10852 8876 10908
rect 8812 10848 8876 10852
rect 8892 10908 8956 10912
rect 8892 10852 8896 10908
rect 8896 10852 8952 10908
rect 8952 10852 8956 10908
rect 8892 10848 8956 10852
rect 8972 10908 9036 10912
rect 8972 10852 8976 10908
rect 8976 10852 9032 10908
rect 9032 10852 9036 10908
rect 8972 10848 9036 10852
rect 14652 10908 14716 10912
rect 14652 10852 14656 10908
rect 14656 10852 14712 10908
rect 14712 10852 14716 10908
rect 14652 10848 14716 10852
rect 14732 10908 14796 10912
rect 14732 10852 14736 10908
rect 14736 10852 14792 10908
rect 14792 10852 14796 10908
rect 14732 10848 14796 10852
rect 14812 10908 14876 10912
rect 14812 10852 14816 10908
rect 14816 10852 14872 10908
rect 14872 10852 14876 10908
rect 14812 10848 14876 10852
rect 14892 10908 14956 10912
rect 14892 10852 14896 10908
rect 14896 10852 14952 10908
rect 14952 10852 14956 10908
rect 14892 10848 14956 10852
rect 14972 10908 15036 10912
rect 14972 10852 14976 10908
rect 14976 10852 15032 10908
rect 15032 10852 15036 10908
rect 14972 10848 15036 10852
rect 1912 10364 1976 10368
rect 1912 10308 1916 10364
rect 1916 10308 1972 10364
rect 1972 10308 1976 10364
rect 1912 10304 1976 10308
rect 1992 10364 2056 10368
rect 1992 10308 1996 10364
rect 1996 10308 2052 10364
rect 2052 10308 2056 10364
rect 1992 10304 2056 10308
rect 2072 10364 2136 10368
rect 2072 10308 2076 10364
rect 2076 10308 2132 10364
rect 2132 10308 2136 10364
rect 2072 10304 2136 10308
rect 2152 10364 2216 10368
rect 2152 10308 2156 10364
rect 2156 10308 2212 10364
rect 2212 10308 2216 10364
rect 2152 10304 2216 10308
rect 2232 10364 2296 10368
rect 2232 10308 2236 10364
rect 2236 10308 2292 10364
rect 2292 10308 2296 10364
rect 2232 10304 2296 10308
rect 7912 10364 7976 10368
rect 7912 10308 7916 10364
rect 7916 10308 7972 10364
rect 7972 10308 7976 10364
rect 7912 10304 7976 10308
rect 7992 10364 8056 10368
rect 7992 10308 7996 10364
rect 7996 10308 8052 10364
rect 8052 10308 8056 10364
rect 7992 10304 8056 10308
rect 8072 10364 8136 10368
rect 8072 10308 8076 10364
rect 8076 10308 8132 10364
rect 8132 10308 8136 10364
rect 8072 10304 8136 10308
rect 8152 10364 8216 10368
rect 8152 10308 8156 10364
rect 8156 10308 8212 10364
rect 8212 10308 8216 10364
rect 8152 10304 8216 10308
rect 8232 10364 8296 10368
rect 8232 10308 8236 10364
rect 8236 10308 8292 10364
rect 8292 10308 8296 10364
rect 8232 10304 8296 10308
rect 13912 10364 13976 10368
rect 13912 10308 13916 10364
rect 13916 10308 13972 10364
rect 13972 10308 13976 10364
rect 13912 10304 13976 10308
rect 13992 10364 14056 10368
rect 13992 10308 13996 10364
rect 13996 10308 14052 10364
rect 14052 10308 14056 10364
rect 13992 10304 14056 10308
rect 14072 10364 14136 10368
rect 14072 10308 14076 10364
rect 14076 10308 14132 10364
rect 14132 10308 14136 10364
rect 14072 10304 14136 10308
rect 14152 10364 14216 10368
rect 14152 10308 14156 10364
rect 14156 10308 14212 10364
rect 14212 10308 14216 10364
rect 14152 10304 14216 10308
rect 14232 10364 14296 10368
rect 14232 10308 14236 10364
rect 14236 10308 14292 10364
rect 14292 10308 14296 10364
rect 14232 10304 14296 10308
rect 2652 9820 2716 9824
rect 2652 9764 2656 9820
rect 2656 9764 2712 9820
rect 2712 9764 2716 9820
rect 2652 9760 2716 9764
rect 2732 9820 2796 9824
rect 2732 9764 2736 9820
rect 2736 9764 2792 9820
rect 2792 9764 2796 9820
rect 2732 9760 2796 9764
rect 2812 9820 2876 9824
rect 2812 9764 2816 9820
rect 2816 9764 2872 9820
rect 2872 9764 2876 9820
rect 2812 9760 2876 9764
rect 2892 9820 2956 9824
rect 2892 9764 2896 9820
rect 2896 9764 2952 9820
rect 2952 9764 2956 9820
rect 2892 9760 2956 9764
rect 2972 9820 3036 9824
rect 2972 9764 2976 9820
rect 2976 9764 3032 9820
rect 3032 9764 3036 9820
rect 2972 9760 3036 9764
rect 8652 9820 8716 9824
rect 8652 9764 8656 9820
rect 8656 9764 8712 9820
rect 8712 9764 8716 9820
rect 8652 9760 8716 9764
rect 8732 9820 8796 9824
rect 8732 9764 8736 9820
rect 8736 9764 8792 9820
rect 8792 9764 8796 9820
rect 8732 9760 8796 9764
rect 8812 9820 8876 9824
rect 8812 9764 8816 9820
rect 8816 9764 8872 9820
rect 8872 9764 8876 9820
rect 8812 9760 8876 9764
rect 8892 9820 8956 9824
rect 8892 9764 8896 9820
rect 8896 9764 8952 9820
rect 8952 9764 8956 9820
rect 8892 9760 8956 9764
rect 8972 9820 9036 9824
rect 8972 9764 8976 9820
rect 8976 9764 9032 9820
rect 9032 9764 9036 9820
rect 8972 9760 9036 9764
rect 14652 9820 14716 9824
rect 14652 9764 14656 9820
rect 14656 9764 14712 9820
rect 14712 9764 14716 9820
rect 14652 9760 14716 9764
rect 14732 9820 14796 9824
rect 14732 9764 14736 9820
rect 14736 9764 14792 9820
rect 14792 9764 14796 9820
rect 14732 9760 14796 9764
rect 14812 9820 14876 9824
rect 14812 9764 14816 9820
rect 14816 9764 14872 9820
rect 14872 9764 14876 9820
rect 14812 9760 14876 9764
rect 14892 9820 14956 9824
rect 14892 9764 14896 9820
rect 14896 9764 14952 9820
rect 14952 9764 14956 9820
rect 14892 9760 14956 9764
rect 14972 9820 15036 9824
rect 14972 9764 14976 9820
rect 14976 9764 15032 9820
rect 15032 9764 15036 9820
rect 14972 9760 15036 9764
rect 14412 9420 14476 9484
rect 1912 9276 1976 9280
rect 1912 9220 1916 9276
rect 1916 9220 1972 9276
rect 1972 9220 1976 9276
rect 1912 9216 1976 9220
rect 1992 9276 2056 9280
rect 1992 9220 1996 9276
rect 1996 9220 2052 9276
rect 2052 9220 2056 9276
rect 1992 9216 2056 9220
rect 2072 9276 2136 9280
rect 2072 9220 2076 9276
rect 2076 9220 2132 9276
rect 2132 9220 2136 9276
rect 2072 9216 2136 9220
rect 2152 9276 2216 9280
rect 2152 9220 2156 9276
rect 2156 9220 2212 9276
rect 2212 9220 2216 9276
rect 2152 9216 2216 9220
rect 2232 9276 2296 9280
rect 2232 9220 2236 9276
rect 2236 9220 2292 9276
rect 2292 9220 2296 9276
rect 2232 9216 2296 9220
rect 7912 9276 7976 9280
rect 7912 9220 7916 9276
rect 7916 9220 7972 9276
rect 7972 9220 7976 9276
rect 7912 9216 7976 9220
rect 7992 9276 8056 9280
rect 7992 9220 7996 9276
rect 7996 9220 8052 9276
rect 8052 9220 8056 9276
rect 7992 9216 8056 9220
rect 8072 9276 8136 9280
rect 8072 9220 8076 9276
rect 8076 9220 8132 9276
rect 8132 9220 8136 9276
rect 8072 9216 8136 9220
rect 8152 9276 8216 9280
rect 8152 9220 8156 9276
rect 8156 9220 8212 9276
rect 8212 9220 8216 9276
rect 8152 9216 8216 9220
rect 8232 9276 8296 9280
rect 8232 9220 8236 9276
rect 8236 9220 8292 9276
rect 8292 9220 8296 9276
rect 8232 9216 8296 9220
rect 13912 9276 13976 9280
rect 13912 9220 13916 9276
rect 13916 9220 13972 9276
rect 13972 9220 13976 9276
rect 13912 9216 13976 9220
rect 13992 9276 14056 9280
rect 13992 9220 13996 9276
rect 13996 9220 14052 9276
rect 14052 9220 14056 9276
rect 13992 9216 14056 9220
rect 14072 9276 14136 9280
rect 14072 9220 14076 9276
rect 14076 9220 14132 9276
rect 14132 9220 14136 9276
rect 14072 9216 14136 9220
rect 14152 9276 14216 9280
rect 14152 9220 14156 9276
rect 14156 9220 14212 9276
rect 14212 9220 14216 9276
rect 14152 9216 14216 9220
rect 14232 9276 14296 9280
rect 14232 9220 14236 9276
rect 14236 9220 14292 9276
rect 14292 9220 14296 9276
rect 14232 9216 14296 9220
rect 2652 8732 2716 8736
rect 2652 8676 2656 8732
rect 2656 8676 2712 8732
rect 2712 8676 2716 8732
rect 2652 8672 2716 8676
rect 2732 8732 2796 8736
rect 2732 8676 2736 8732
rect 2736 8676 2792 8732
rect 2792 8676 2796 8732
rect 2732 8672 2796 8676
rect 2812 8732 2876 8736
rect 2812 8676 2816 8732
rect 2816 8676 2872 8732
rect 2872 8676 2876 8732
rect 2812 8672 2876 8676
rect 2892 8732 2956 8736
rect 2892 8676 2896 8732
rect 2896 8676 2952 8732
rect 2952 8676 2956 8732
rect 2892 8672 2956 8676
rect 2972 8732 3036 8736
rect 2972 8676 2976 8732
rect 2976 8676 3032 8732
rect 3032 8676 3036 8732
rect 2972 8672 3036 8676
rect 8652 8732 8716 8736
rect 8652 8676 8656 8732
rect 8656 8676 8712 8732
rect 8712 8676 8716 8732
rect 8652 8672 8716 8676
rect 8732 8732 8796 8736
rect 8732 8676 8736 8732
rect 8736 8676 8792 8732
rect 8792 8676 8796 8732
rect 8732 8672 8796 8676
rect 8812 8732 8876 8736
rect 8812 8676 8816 8732
rect 8816 8676 8872 8732
rect 8872 8676 8876 8732
rect 8812 8672 8876 8676
rect 8892 8732 8956 8736
rect 8892 8676 8896 8732
rect 8896 8676 8952 8732
rect 8952 8676 8956 8732
rect 8892 8672 8956 8676
rect 8972 8732 9036 8736
rect 8972 8676 8976 8732
rect 8976 8676 9032 8732
rect 9032 8676 9036 8732
rect 8972 8672 9036 8676
rect 14652 8732 14716 8736
rect 14652 8676 14656 8732
rect 14656 8676 14712 8732
rect 14712 8676 14716 8732
rect 14652 8672 14716 8676
rect 14732 8732 14796 8736
rect 14732 8676 14736 8732
rect 14736 8676 14792 8732
rect 14792 8676 14796 8732
rect 14732 8672 14796 8676
rect 14812 8732 14876 8736
rect 14812 8676 14816 8732
rect 14816 8676 14872 8732
rect 14872 8676 14876 8732
rect 14812 8672 14876 8676
rect 14892 8732 14956 8736
rect 14892 8676 14896 8732
rect 14896 8676 14952 8732
rect 14952 8676 14956 8732
rect 14892 8672 14956 8676
rect 14972 8732 15036 8736
rect 14972 8676 14976 8732
rect 14976 8676 15032 8732
rect 15032 8676 15036 8732
rect 14972 8672 15036 8676
rect 1912 8188 1976 8192
rect 1912 8132 1916 8188
rect 1916 8132 1972 8188
rect 1972 8132 1976 8188
rect 1912 8128 1976 8132
rect 1992 8188 2056 8192
rect 1992 8132 1996 8188
rect 1996 8132 2052 8188
rect 2052 8132 2056 8188
rect 1992 8128 2056 8132
rect 2072 8188 2136 8192
rect 2072 8132 2076 8188
rect 2076 8132 2132 8188
rect 2132 8132 2136 8188
rect 2072 8128 2136 8132
rect 2152 8188 2216 8192
rect 2152 8132 2156 8188
rect 2156 8132 2212 8188
rect 2212 8132 2216 8188
rect 2152 8128 2216 8132
rect 2232 8188 2296 8192
rect 2232 8132 2236 8188
rect 2236 8132 2292 8188
rect 2292 8132 2296 8188
rect 2232 8128 2296 8132
rect 7912 8188 7976 8192
rect 7912 8132 7916 8188
rect 7916 8132 7972 8188
rect 7972 8132 7976 8188
rect 7912 8128 7976 8132
rect 7992 8188 8056 8192
rect 7992 8132 7996 8188
rect 7996 8132 8052 8188
rect 8052 8132 8056 8188
rect 7992 8128 8056 8132
rect 8072 8188 8136 8192
rect 8072 8132 8076 8188
rect 8076 8132 8132 8188
rect 8132 8132 8136 8188
rect 8072 8128 8136 8132
rect 8152 8188 8216 8192
rect 8152 8132 8156 8188
rect 8156 8132 8212 8188
rect 8212 8132 8216 8188
rect 8152 8128 8216 8132
rect 8232 8188 8296 8192
rect 8232 8132 8236 8188
rect 8236 8132 8292 8188
rect 8292 8132 8296 8188
rect 8232 8128 8296 8132
rect 13912 8188 13976 8192
rect 13912 8132 13916 8188
rect 13916 8132 13972 8188
rect 13972 8132 13976 8188
rect 13912 8128 13976 8132
rect 13992 8188 14056 8192
rect 13992 8132 13996 8188
rect 13996 8132 14052 8188
rect 14052 8132 14056 8188
rect 13992 8128 14056 8132
rect 14072 8188 14136 8192
rect 14072 8132 14076 8188
rect 14076 8132 14132 8188
rect 14132 8132 14136 8188
rect 14072 8128 14136 8132
rect 14152 8188 14216 8192
rect 14152 8132 14156 8188
rect 14156 8132 14212 8188
rect 14212 8132 14216 8188
rect 14152 8128 14216 8132
rect 14232 8188 14296 8192
rect 14232 8132 14236 8188
rect 14236 8132 14292 8188
rect 14292 8132 14296 8188
rect 14232 8128 14296 8132
rect 12572 7652 12636 7716
rect 2652 7644 2716 7648
rect 2652 7588 2656 7644
rect 2656 7588 2712 7644
rect 2712 7588 2716 7644
rect 2652 7584 2716 7588
rect 2732 7644 2796 7648
rect 2732 7588 2736 7644
rect 2736 7588 2792 7644
rect 2792 7588 2796 7644
rect 2732 7584 2796 7588
rect 2812 7644 2876 7648
rect 2812 7588 2816 7644
rect 2816 7588 2872 7644
rect 2872 7588 2876 7644
rect 2812 7584 2876 7588
rect 2892 7644 2956 7648
rect 2892 7588 2896 7644
rect 2896 7588 2952 7644
rect 2952 7588 2956 7644
rect 2892 7584 2956 7588
rect 2972 7644 3036 7648
rect 2972 7588 2976 7644
rect 2976 7588 3032 7644
rect 3032 7588 3036 7644
rect 2972 7584 3036 7588
rect 8652 7644 8716 7648
rect 8652 7588 8656 7644
rect 8656 7588 8712 7644
rect 8712 7588 8716 7644
rect 8652 7584 8716 7588
rect 8732 7644 8796 7648
rect 8732 7588 8736 7644
rect 8736 7588 8792 7644
rect 8792 7588 8796 7644
rect 8732 7584 8796 7588
rect 8812 7644 8876 7648
rect 8812 7588 8816 7644
rect 8816 7588 8872 7644
rect 8872 7588 8876 7644
rect 8812 7584 8876 7588
rect 8892 7644 8956 7648
rect 8892 7588 8896 7644
rect 8896 7588 8952 7644
rect 8952 7588 8956 7644
rect 8892 7584 8956 7588
rect 8972 7644 9036 7648
rect 8972 7588 8976 7644
rect 8976 7588 9032 7644
rect 9032 7588 9036 7644
rect 8972 7584 9036 7588
rect 14652 7644 14716 7648
rect 14652 7588 14656 7644
rect 14656 7588 14712 7644
rect 14712 7588 14716 7644
rect 14652 7584 14716 7588
rect 14732 7644 14796 7648
rect 14732 7588 14736 7644
rect 14736 7588 14792 7644
rect 14792 7588 14796 7644
rect 14732 7584 14796 7588
rect 14812 7644 14876 7648
rect 14812 7588 14816 7644
rect 14816 7588 14872 7644
rect 14872 7588 14876 7644
rect 14812 7584 14876 7588
rect 14892 7644 14956 7648
rect 14892 7588 14896 7644
rect 14896 7588 14952 7644
rect 14952 7588 14956 7644
rect 14892 7584 14956 7588
rect 14972 7644 15036 7648
rect 14972 7588 14976 7644
rect 14976 7588 15032 7644
rect 15032 7588 15036 7644
rect 14972 7584 15036 7588
rect 1912 7100 1976 7104
rect 1912 7044 1916 7100
rect 1916 7044 1972 7100
rect 1972 7044 1976 7100
rect 1912 7040 1976 7044
rect 1992 7100 2056 7104
rect 1992 7044 1996 7100
rect 1996 7044 2052 7100
rect 2052 7044 2056 7100
rect 1992 7040 2056 7044
rect 2072 7100 2136 7104
rect 2072 7044 2076 7100
rect 2076 7044 2132 7100
rect 2132 7044 2136 7100
rect 2072 7040 2136 7044
rect 2152 7100 2216 7104
rect 2152 7044 2156 7100
rect 2156 7044 2212 7100
rect 2212 7044 2216 7100
rect 2152 7040 2216 7044
rect 2232 7100 2296 7104
rect 2232 7044 2236 7100
rect 2236 7044 2292 7100
rect 2292 7044 2296 7100
rect 2232 7040 2296 7044
rect 7912 7100 7976 7104
rect 7912 7044 7916 7100
rect 7916 7044 7972 7100
rect 7972 7044 7976 7100
rect 7912 7040 7976 7044
rect 7992 7100 8056 7104
rect 7992 7044 7996 7100
rect 7996 7044 8052 7100
rect 8052 7044 8056 7100
rect 7992 7040 8056 7044
rect 8072 7100 8136 7104
rect 8072 7044 8076 7100
rect 8076 7044 8132 7100
rect 8132 7044 8136 7100
rect 8072 7040 8136 7044
rect 8152 7100 8216 7104
rect 8152 7044 8156 7100
rect 8156 7044 8212 7100
rect 8212 7044 8216 7100
rect 8152 7040 8216 7044
rect 8232 7100 8296 7104
rect 8232 7044 8236 7100
rect 8236 7044 8292 7100
rect 8292 7044 8296 7100
rect 8232 7040 8296 7044
rect 13912 7100 13976 7104
rect 13912 7044 13916 7100
rect 13916 7044 13972 7100
rect 13972 7044 13976 7100
rect 13912 7040 13976 7044
rect 13992 7100 14056 7104
rect 13992 7044 13996 7100
rect 13996 7044 14052 7100
rect 14052 7044 14056 7100
rect 13992 7040 14056 7044
rect 14072 7100 14136 7104
rect 14072 7044 14076 7100
rect 14076 7044 14132 7100
rect 14132 7044 14136 7100
rect 14072 7040 14136 7044
rect 14152 7100 14216 7104
rect 14152 7044 14156 7100
rect 14156 7044 14212 7100
rect 14212 7044 14216 7100
rect 14152 7040 14216 7044
rect 14232 7100 14296 7104
rect 14232 7044 14236 7100
rect 14236 7044 14292 7100
rect 14292 7044 14296 7100
rect 14232 7040 14296 7044
rect 2652 6556 2716 6560
rect 2652 6500 2656 6556
rect 2656 6500 2712 6556
rect 2712 6500 2716 6556
rect 2652 6496 2716 6500
rect 2732 6556 2796 6560
rect 2732 6500 2736 6556
rect 2736 6500 2792 6556
rect 2792 6500 2796 6556
rect 2732 6496 2796 6500
rect 2812 6556 2876 6560
rect 2812 6500 2816 6556
rect 2816 6500 2872 6556
rect 2872 6500 2876 6556
rect 2812 6496 2876 6500
rect 2892 6556 2956 6560
rect 2892 6500 2896 6556
rect 2896 6500 2952 6556
rect 2952 6500 2956 6556
rect 2892 6496 2956 6500
rect 2972 6556 3036 6560
rect 2972 6500 2976 6556
rect 2976 6500 3032 6556
rect 3032 6500 3036 6556
rect 2972 6496 3036 6500
rect 8652 6556 8716 6560
rect 8652 6500 8656 6556
rect 8656 6500 8712 6556
rect 8712 6500 8716 6556
rect 8652 6496 8716 6500
rect 8732 6556 8796 6560
rect 8732 6500 8736 6556
rect 8736 6500 8792 6556
rect 8792 6500 8796 6556
rect 8732 6496 8796 6500
rect 8812 6556 8876 6560
rect 8812 6500 8816 6556
rect 8816 6500 8872 6556
rect 8872 6500 8876 6556
rect 8812 6496 8876 6500
rect 8892 6556 8956 6560
rect 8892 6500 8896 6556
rect 8896 6500 8952 6556
rect 8952 6500 8956 6556
rect 8892 6496 8956 6500
rect 8972 6556 9036 6560
rect 8972 6500 8976 6556
rect 8976 6500 9032 6556
rect 9032 6500 9036 6556
rect 8972 6496 9036 6500
rect 14652 6556 14716 6560
rect 14652 6500 14656 6556
rect 14656 6500 14712 6556
rect 14712 6500 14716 6556
rect 14652 6496 14716 6500
rect 14732 6556 14796 6560
rect 14732 6500 14736 6556
rect 14736 6500 14792 6556
rect 14792 6500 14796 6556
rect 14732 6496 14796 6500
rect 14812 6556 14876 6560
rect 14812 6500 14816 6556
rect 14816 6500 14872 6556
rect 14872 6500 14876 6556
rect 14812 6496 14876 6500
rect 14892 6556 14956 6560
rect 14892 6500 14896 6556
rect 14896 6500 14952 6556
rect 14952 6500 14956 6556
rect 14892 6496 14956 6500
rect 14972 6556 15036 6560
rect 14972 6500 14976 6556
rect 14976 6500 15032 6556
rect 15032 6500 15036 6556
rect 14972 6496 15036 6500
rect 14412 6488 14476 6492
rect 14412 6432 14462 6488
rect 14462 6432 14476 6488
rect 14412 6428 14476 6432
rect 1912 6012 1976 6016
rect 1912 5956 1916 6012
rect 1916 5956 1972 6012
rect 1972 5956 1976 6012
rect 1912 5952 1976 5956
rect 1992 6012 2056 6016
rect 1992 5956 1996 6012
rect 1996 5956 2052 6012
rect 2052 5956 2056 6012
rect 1992 5952 2056 5956
rect 2072 6012 2136 6016
rect 2072 5956 2076 6012
rect 2076 5956 2132 6012
rect 2132 5956 2136 6012
rect 2072 5952 2136 5956
rect 2152 6012 2216 6016
rect 2152 5956 2156 6012
rect 2156 5956 2212 6012
rect 2212 5956 2216 6012
rect 2152 5952 2216 5956
rect 2232 6012 2296 6016
rect 2232 5956 2236 6012
rect 2236 5956 2292 6012
rect 2292 5956 2296 6012
rect 2232 5952 2296 5956
rect 7912 6012 7976 6016
rect 7912 5956 7916 6012
rect 7916 5956 7972 6012
rect 7972 5956 7976 6012
rect 7912 5952 7976 5956
rect 7992 6012 8056 6016
rect 7992 5956 7996 6012
rect 7996 5956 8052 6012
rect 8052 5956 8056 6012
rect 7992 5952 8056 5956
rect 8072 6012 8136 6016
rect 8072 5956 8076 6012
rect 8076 5956 8132 6012
rect 8132 5956 8136 6012
rect 8072 5952 8136 5956
rect 8152 6012 8216 6016
rect 8152 5956 8156 6012
rect 8156 5956 8212 6012
rect 8212 5956 8216 6012
rect 8152 5952 8216 5956
rect 8232 6012 8296 6016
rect 8232 5956 8236 6012
rect 8236 5956 8292 6012
rect 8292 5956 8296 6012
rect 8232 5952 8296 5956
rect 13912 6012 13976 6016
rect 13912 5956 13916 6012
rect 13916 5956 13972 6012
rect 13972 5956 13976 6012
rect 13912 5952 13976 5956
rect 13992 6012 14056 6016
rect 13992 5956 13996 6012
rect 13996 5956 14052 6012
rect 14052 5956 14056 6012
rect 13992 5952 14056 5956
rect 14072 6012 14136 6016
rect 14072 5956 14076 6012
rect 14076 5956 14132 6012
rect 14132 5956 14136 6012
rect 14072 5952 14136 5956
rect 14152 6012 14216 6016
rect 14152 5956 14156 6012
rect 14156 5956 14212 6012
rect 14212 5956 14216 6012
rect 14152 5952 14216 5956
rect 14232 6012 14296 6016
rect 14232 5956 14236 6012
rect 14236 5956 14292 6012
rect 14292 5956 14296 6012
rect 14232 5952 14296 5956
rect 2652 5468 2716 5472
rect 2652 5412 2656 5468
rect 2656 5412 2712 5468
rect 2712 5412 2716 5468
rect 2652 5408 2716 5412
rect 2732 5468 2796 5472
rect 2732 5412 2736 5468
rect 2736 5412 2792 5468
rect 2792 5412 2796 5468
rect 2732 5408 2796 5412
rect 2812 5468 2876 5472
rect 2812 5412 2816 5468
rect 2816 5412 2872 5468
rect 2872 5412 2876 5468
rect 2812 5408 2876 5412
rect 2892 5468 2956 5472
rect 2892 5412 2896 5468
rect 2896 5412 2952 5468
rect 2952 5412 2956 5468
rect 2892 5408 2956 5412
rect 2972 5468 3036 5472
rect 2972 5412 2976 5468
rect 2976 5412 3032 5468
rect 3032 5412 3036 5468
rect 2972 5408 3036 5412
rect 8652 5468 8716 5472
rect 8652 5412 8656 5468
rect 8656 5412 8712 5468
rect 8712 5412 8716 5468
rect 8652 5408 8716 5412
rect 8732 5468 8796 5472
rect 8732 5412 8736 5468
rect 8736 5412 8792 5468
rect 8792 5412 8796 5468
rect 8732 5408 8796 5412
rect 8812 5468 8876 5472
rect 8812 5412 8816 5468
rect 8816 5412 8872 5468
rect 8872 5412 8876 5468
rect 8812 5408 8876 5412
rect 8892 5468 8956 5472
rect 8892 5412 8896 5468
rect 8896 5412 8952 5468
rect 8952 5412 8956 5468
rect 8892 5408 8956 5412
rect 8972 5468 9036 5472
rect 8972 5412 8976 5468
rect 8976 5412 9032 5468
rect 9032 5412 9036 5468
rect 8972 5408 9036 5412
rect 14652 5468 14716 5472
rect 14652 5412 14656 5468
rect 14656 5412 14712 5468
rect 14712 5412 14716 5468
rect 14652 5408 14716 5412
rect 14732 5468 14796 5472
rect 14732 5412 14736 5468
rect 14736 5412 14792 5468
rect 14792 5412 14796 5468
rect 14732 5408 14796 5412
rect 14812 5468 14876 5472
rect 14812 5412 14816 5468
rect 14816 5412 14872 5468
rect 14872 5412 14876 5468
rect 14812 5408 14876 5412
rect 14892 5468 14956 5472
rect 14892 5412 14896 5468
rect 14896 5412 14952 5468
rect 14952 5412 14956 5468
rect 14892 5408 14956 5412
rect 14972 5468 15036 5472
rect 14972 5412 14976 5468
rect 14976 5412 15032 5468
rect 15032 5412 15036 5468
rect 14972 5408 15036 5412
rect 1912 4924 1976 4928
rect 1912 4868 1916 4924
rect 1916 4868 1972 4924
rect 1972 4868 1976 4924
rect 1912 4864 1976 4868
rect 1992 4924 2056 4928
rect 1992 4868 1996 4924
rect 1996 4868 2052 4924
rect 2052 4868 2056 4924
rect 1992 4864 2056 4868
rect 2072 4924 2136 4928
rect 2072 4868 2076 4924
rect 2076 4868 2132 4924
rect 2132 4868 2136 4924
rect 2072 4864 2136 4868
rect 2152 4924 2216 4928
rect 2152 4868 2156 4924
rect 2156 4868 2212 4924
rect 2212 4868 2216 4924
rect 2152 4864 2216 4868
rect 2232 4924 2296 4928
rect 2232 4868 2236 4924
rect 2236 4868 2292 4924
rect 2292 4868 2296 4924
rect 2232 4864 2296 4868
rect 7912 4924 7976 4928
rect 7912 4868 7916 4924
rect 7916 4868 7972 4924
rect 7972 4868 7976 4924
rect 7912 4864 7976 4868
rect 7992 4924 8056 4928
rect 7992 4868 7996 4924
rect 7996 4868 8052 4924
rect 8052 4868 8056 4924
rect 7992 4864 8056 4868
rect 8072 4924 8136 4928
rect 8072 4868 8076 4924
rect 8076 4868 8132 4924
rect 8132 4868 8136 4924
rect 8072 4864 8136 4868
rect 8152 4924 8216 4928
rect 8152 4868 8156 4924
rect 8156 4868 8212 4924
rect 8212 4868 8216 4924
rect 8152 4864 8216 4868
rect 8232 4924 8296 4928
rect 8232 4868 8236 4924
rect 8236 4868 8292 4924
rect 8292 4868 8296 4924
rect 8232 4864 8296 4868
rect 13912 4924 13976 4928
rect 13912 4868 13916 4924
rect 13916 4868 13972 4924
rect 13972 4868 13976 4924
rect 13912 4864 13976 4868
rect 13992 4924 14056 4928
rect 13992 4868 13996 4924
rect 13996 4868 14052 4924
rect 14052 4868 14056 4924
rect 13992 4864 14056 4868
rect 14072 4924 14136 4928
rect 14072 4868 14076 4924
rect 14076 4868 14132 4924
rect 14132 4868 14136 4924
rect 14072 4864 14136 4868
rect 14152 4924 14216 4928
rect 14152 4868 14156 4924
rect 14156 4868 14212 4924
rect 14212 4868 14216 4924
rect 14152 4864 14216 4868
rect 14232 4924 14296 4928
rect 14232 4868 14236 4924
rect 14236 4868 14292 4924
rect 14292 4868 14296 4924
rect 14232 4864 14296 4868
rect 2652 4380 2716 4384
rect 2652 4324 2656 4380
rect 2656 4324 2712 4380
rect 2712 4324 2716 4380
rect 2652 4320 2716 4324
rect 2732 4380 2796 4384
rect 2732 4324 2736 4380
rect 2736 4324 2792 4380
rect 2792 4324 2796 4380
rect 2732 4320 2796 4324
rect 2812 4380 2876 4384
rect 2812 4324 2816 4380
rect 2816 4324 2872 4380
rect 2872 4324 2876 4380
rect 2812 4320 2876 4324
rect 2892 4380 2956 4384
rect 2892 4324 2896 4380
rect 2896 4324 2952 4380
rect 2952 4324 2956 4380
rect 2892 4320 2956 4324
rect 2972 4380 3036 4384
rect 2972 4324 2976 4380
rect 2976 4324 3032 4380
rect 3032 4324 3036 4380
rect 2972 4320 3036 4324
rect 8652 4380 8716 4384
rect 8652 4324 8656 4380
rect 8656 4324 8712 4380
rect 8712 4324 8716 4380
rect 8652 4320 8716 4324
rect 8732 4380 8796 4384
rect 8732 4324 8736 4380
rect 8736 4324 8792 4380
rect 8792 4324 8796 4380
rect 8732 4320 8796 4324
rect 8812 4380 8876 4384
rect 8812 4324 8816 4380
rect 8816 4324 8872 4380
rect 8872 4324 8876 4380
rect 8812 4320 8876 4324
rect 8892 4380 8956 4384
rect 8892 4324 8896 4380
rect 8896 4324 8952 4380
rect 8952 4324 8956 4380
rect 8892 4320 8956 4324
rect 8972 4380 9036 4384
rect 8972 4324 8976 4380
rect 8976 4324 9032 4380
rect 9032 4324 9036 4380
rect 8972 4320 9036 4324
rect 14652 4380 14716 4384
rect 14652 4324 14656 4380
rect 14656 4324 14712 4380
rect 14712 4324 14716 4380
rect 14652 4320 14716 4324
rect 14732 4380 14796 4384
rect 14732 4324 14736 4380
rect 14736 4324 14792 4380
rect 14792 4324 14796 4380
rect 14732 4320 14796 4324
rect 14812 4380 14876 4384
rect 14812 4324 14816 4380
rect 14816 4324 14872 4380
rect 14872 4324 14876 4380
rect 14812 4320 14876 4324
rect 14892 4380 14956 4384
rect 14892 4324 14896 4380
rect 14896 4324 14952 4380
rect 14952 4324 14956 4380
rect 14892 4320 14956 4324
rect 14972 4380 15036 4384
rect 14972 4324 14976 4380
rect 14976 4324 15032 4380
rect 15032 4324 15036 4380
rect 14972 4320 15036 4324
rect 1912 3836 1976 3840
rect 1912 3780 1916 3836
rect 1916 3780 1972 3836
rect 1972 3780 1976 3836
rect 1912 3776 1976 3780
rect 1992 3836 2056 3840
rect 1992 3780 1996 3836
rect 1996 3780 2052 3836
rect 2052 3780 2056 3836
rect 1992 3776 2056 3780
rect 2072 3836 2136 3840
rect 2072 3780 2076 3836
rect 2076 3780 2132 3836
rect 2132 3780 2136 3836
rect 2072 3776 2136 3780
rect 2152 3836 2216 3840
rect 2152 3780 2156 3836
rect 2156 3780 2212 3836
rect 2212 3780 2216 3836
rect 2152 3776 2216 3780
rect 2232 3836 2296 3840
rect 2232 3780 2236 3836
rect 2236 3780 2292 3836
rect 2292 3780 2296 3836
rect 2232 3776 2296 3780
rect 7912 3836 7976 3840
rect 7912 3780 7916 3836
rect 7916 3780 7972 3836
rect 7972 3780 7976 3836
rect 7912 3776 7976 3780
rect 7992 3836 8056 3840
rect 7992 3780 7996 3836
rect 7996 3780 8052 3836
rect 8052 3780 8056 3836
rect 7992 3776 8056 3780
rect 8072 3836 8136 3840
rect 8072 3780 8076 3836
rect 8076 3780 8132 3836
rect 8132 3780 8136 3836
rect 8072 3776 8136 3780
rect 8152 3836 8216 3840
rect 8152 3780 8156 3836
rect 8156 3780 8212 3836
rect 8212 3780 8216 3836
rect 8152 3776 8216 3780
rect 8232 3836 8296 3840
rect 8232 3780 8236 3836
rect 8236 3780 8292 3836
rect 8292 3780 8296 3836
rect 8232 3776 8296 3780
rect 13912 3836 13976 3840
rect 13912 3780 13916 3836
rect 13916 3780 13972 3836
rect 13972 3780 13976 3836
rect 13912 3776 13976 3780
rect 13992 3836 14056 3840
rect 13992 3780 13996 3836
rect 13996 3780 14052 3836
rect 14052 3780 14056 3836
rect 13992 3776 14056 3780
rect 14072 3836 14136 3840
rect 14072 3780 14076 3836
rect 14076 3780 14132 3836
rect 14132 3780 14136 3836
rect 14072 3776 14136 3780
rect 14152 3836 14216 3840
rect 14152 3780 14156 3836
rect 14156 3780 14212 3836
rect 14212 3780 14216 3836
rect 14152 3776 14216 3780
rect 14232 3836 14296 3840
rect 14232 3780 14236 3836
rect 14236 3780 14292 3836
rect 14292 3780 14296 3836
rect 14232 3776 14296 3780
rect 2652 3292 2716 3296
rect 2652 3236 2656 3292
rect 2656 3236 2712 3292
rect 2712 3236 2716 3292
rect 2652 3232 2716 3236
rect 2732 3292 2796 3296
rect 2732 3236 2736 3292
rect 2736 3236 2792 3292
rect 2792 3236 2796 3292
rect 2732 3232 2796 3236
rect 2812 3292 2876 3296
rect 2812 3236 2816 3292
rect 2816 3236 2872 3292
rect 2872 3236 2876 3292
rect 2812 3232 2876 3236
rect 2892 3292 2956 3296
rect 2892 3236 2896 3292
rect 2896 3236 2952 3292
rect 2952 3236 2956 3292
rect 2892 3232 2956 3236
rect 2972 3292 3036 3296
rect 2972 3236 2976 3292
rect 2976 3236 3032 3292
rect 3032 3236 3036 3292
rect 2972 3232 3036 3236
rect 8652 3292 8716 3296
rect 8652 3236 8656 3292
rect 8656 3236 8712 3292
rect 8712 3236 8716 3292
rect 8652 3232 8716 3236
rect 8732 3292 8796 3296
rect 8732 3236 8736 3292
rect 8736 3236 8792 3292
rect 8792 3236 8796 3292
rect 8732 3232 8796 3236
rect 8812 3292 8876 3296
rect 8812 3236 8816 3292
rect 8816 3236 8872 3292
rect 8872 3236 8876 3292
rect 8812 3232 8876 3236
rect 8892 3292 8956 3296
rect 8892 3236 8896 3292
rect 8896 3236 8952 3292
rect 8952 3236 8956 3292
rect 8892 3232 8956 3236
rect 8972 3292 9036 3296
rect 8972 3236 8976 3292
rect 8976 3236 9032 3292
rect 9032 3236 9036 3292
rect 8972 3232 9036 3236
rect 14652 3292 14716 3296
rect 14652 3236 14656 3292
rect 14656 3236 14712 3292
rect 14712 3236 14716 3292
rect 14652 3232 14716 3236
rect 14732 3292 14796 3296
rect 14732 3236 14736 3292
rect 14736 3236 14792 3292
rect 14792 3236 14796 3292
rect 14732 3232 14796 3236
rect 14812 3292 14876 3296
rect 14812 3236 14816 3292
rect 14816 3236 14872 3292
rect 14872 3236 14876 3292
rect 14812 3232 14876 3236
rect 14892 3292 14956 3296
rect 14892 3236 14896 3292
rect 14896 3236 14952 3292
rect 14952 3236 14956 3292
rect 14892 3232 14956 3236
rect 14972 3292 15036 3296
rect 14972 3236 14976 3292
rect 14976 3236 15032 3292
rect 15032 3236 15036 3292
rect 14972 3232 15036 3236
rect 1912 2748 1976 2752
rect 1912 2692 1916 2748
rect 1916 2692 1972 2748
rect 1972 2692 1976 2748
rect 1912 2688 1976 2692
rect 1992 2748 2056 2752
rect 1992 2692 1996 2748
rect 1996 2692 2052 2748
rect 2052 2692 2056 2748
rect 1992 2688 2056 2692
rect 2072 2748 2136 2752
rect 2072 2692 2076 2748
rect 2076 2692 2132 2748
rect 2132 2692 2136 2748
rect 2072 2688 2136 2692
rect 2152 2748 2216 2752
rect 2152 2692 2156 2748
rect 2156 2692 2212 2748
rect 2212 2692 2216 2748
rect 2152 2688 2216 2692
rect 2232 2748 2296 2752
rect 2232 2692 2236 2748
rect 2236 2692 2292 2748
rect 2292 2692 2296 2748
rect 2232 2688 2296 2692
rect 7912 2748 7976 2752
rect 7912 2692 7916 2748
rect 7916 2692 7972 2748
rect 7972 2692 7976 2748
rect 7912 2688 7976 2692
rect 7992 2748 8056 2752
rect 7992 2692 7996 2748
rect 7996 2692 8052 2748
rect 8052 2692 8056 2748
rect 7992 2688 8056 2692
rect 8072 2748 8136 2752
rect 8072 2692 8076 2748
rect 8076 2692 8132 2748
rect 8132 2692 8136 2748
rect 8072 2688 8136 2692
rect 8152 2748 8216 2752
rect 8152 2692 8156 2748
rect 8156 2692 8212 2748
rect 8212 2692 8216 2748
rect 8152 2688 8216 2692
rect 8232 2748 8296 2752
rect 8232 2692 8236 2748
rect 8236 2692 8292 2748
rect 8292 2692 8296 2748
rect 8232 2688 8296 2692
rect 13912 2748 13976 2752
rect 13912 2692 13916 2748
rect 13916 2692 13972 2748
rect 13972 2692 13976 2748
rect 13912 2688 13976 2692
rect 13992 2748 14056 2752
rect 13992 2692 13996 2748
rect 13996 2692 14052 2748
rect 14052 2692 14056 2748
rect 13992 2688 14056 2692
rect 14072 2748 14136 2752
rect 14072 2692 14076 2748
rect 14076 2692 14132 2748
rect 14132 2692 14136 2748
rect 14072 2688 14136 2692
rect 14152 2748 14216 2752
rect 14152 2692 14156 2748
rect 14156 2692 14212 2748
rect 14212 2692 14216 2748
rect 14152 2688 14216 2692
rect 14232 2748 14296 2752
rect 14232 2692 14236 2748
rect 14236 2692 14292 2748
rect 14292 2692 14296 2748
rect 14232 2688 14296 2692
rect 2652 2204 2716 2208
rect 2652 2148 2656 2204
rect 2656 2148 2712 2204
rect 2712 2148 2716 2204
rect 2652 2144 2716 2148
rect 2732 2204 2796 2208
rect 2732 2148 2736 2204
rect 2736 2148 2792 2204
rect 2792 2148 2796 2204
rect 2732 2144 2796 2148
rect 2812 2204 2876 2208
rect 2812 2148 2816 2204
rect 2816 2148 2872 2204
rect 2872 2148 2876 2204
rect 2812 2144 2876 2148
rect 2892 2204 2956 2208
rect 2892 2148 2896 2204
rect 2896 2148 2952 2204
rect 2952 2148 2956 2204
rect 2892 2144 2956 2148
rect 2972 2204 3036 2208
rect 2972 2148 2976 2204
rect 2976 2148 3032 2204
rect 3032 2148 3036 2204
rect 2972 2144 3036 2148
rect 8652 2204 8716 2208
rect 8652 2148 8656 2204
rect 8656 2148 8712 2204
rect 8712 2148 8716 2204
rect 8652 2144 8716 2148
rect 8732 2204 8796 2208
rect 8732 2148 8736 2204
rect 8736 2148 8792 2204
rect 8792 2148 8796 2204
rect 8732 2144 8796 2148
rect 8812 2204 8876 2208
rect 8812 2148 8816 2204
rect 8816 2148 8872 2204
rect 8872 2148 8876 2204
rect 8812 2144 8876 2148
rect 8892 2204 8956 2208
rect 8892 2148 8896 2204
rect 8896 2148 8952 2204
rect 8952 2148 8956 2204
rect 8892 2144 8956 2148
rect 8972 2204 9036 2208
rect 8972 2148 8976 2204
rect 8976 2148 9032 2204
rect 9032 2148 9036 2204
rect 8972 2144 9036 2148
rect 14652 2204 14716 2208
rect 14652 2148 14656 2204
rect 14656 2148 14712 2204
rect 14712 2148 14716 2204
rect 14652 2144 14716 2148
rect 14732 2204 14796 2208
rect 14732 2148 14736 2204
rect 14736 2148 14792 2204
rect 14792 2148 14796 2204
rect 14732 2144 14796 2148
rect 14812 2204 14876 2208
rect 14812 2148 14816 2204
rect 14816 2148 14872 2204
rect 14872 2148 14876 2204
rect 14812 2144 14876 2148
rect 14892 2204 14956 2208
rect 14892 2148 14896 2204
rect 14896 2148 14952 2204
rect 14952 2148 14956 2204
rect 14892 2144 14956 2148
rect 14972 2204 15036 2208
rect 14972 2148 14976 2204
rect 14976 2148 15032 2204
rect 15032 2148 15036 2204
rect 14972 2144 15036 2148
<< metal4 >>
rect 1904 17984 2304 18544
rect 1904 17920 1912 17984
rect 1976 17920 1992 17984
rect 2056 17920 2072 17984
rect 2136 17920 2152 17984
rect 2216 17920 2232 17984
rect 2296 17920 2304 17984
rect 1904 16896 2304 17920
rect 1904 16832 1912 16896
rect 1976 16832 1992 16896
rect 2056 16832 2072 16896
rect 2136 16832 2152 16896
rect 2216 16832 2232 16896
rect 2296 16832 2304 16896
rect 1904 15808 2304 16832
rect 1904 15744 1912 15808
rect 1976 15744 1992 15808
rect 2056 15744 2072 15808
rect 2136 15744 2152 15808
rect 2216 15744 2232 15808
rect 2296 15744 2304 15808
rect 1904 15294 2304 15744
rect 1904 15058 1986 15294
rect 2222 15058 2304 15294
rect 1904 14720 2304 15058
rect 1904 14656 1912 14720
rect 1976 14656 1992 14720
rect 2056 14656 2072 14720
rect 2136 14656 2152 14720
rect 2216 14656 2232 14720
rect 2296 14656 2304 14720
rect 1904 13632 2304 14656
rect 1904 13568 1912 13632
rect 1976 13568 1992 13632
rect 2056 13568 2072 13632
rect 2136 13568 2152 13632
rect 2216 13568 2232 13632
rect 2296 13568 2304 13632
rect 1904 12544 2304 13568
rect 1904 12480 1912 12544
rect 1976 12480 1992 12544
rect 2056 12480 2072 12544
rect 2136 12480 2152 12544
rect 2216 12480 2232 12544
rect 2296 12480 2304 12544
rect 1904 11456 2304 12480
rect 1904 11392 1912 11456
rect 1976 11392 1992 11456
rect 2056 11392 2072 11456
rect 2136 11392 2152 11456
rect 2216 11392 2232 11456
rect 2296 11392 2304 11456
rect 1904 10368 2304 11392
rect 1904 10304 1912 10368
rect 1976 10304 1992 10368
rect 2056 10304 2072 10368
rect 2136 10304 2152 10368
rect 2216 10304 2232 10368
rect 2296 10304 2304 10368
rect 1904 9294 2304 10304
rect 1904 9280 1986 9294
rect 2222 9280 2304 9294
rect 1904 9216 1912 9280
rect 1976 9216 1986 9280
rect 2222 9216 2232 9280
rect 2296 9216 2304 9280
rect 1904 9058 1986 9216
rect 2222 9058 2304 9216
rect 1904 8192 2304 9058
rect 1904 8128 1912 8192
rect 1976 8128 1992 8192
rect 2056 8128 2072 8192
rect 2136 8128 2152 8192
rect 2216 8128 2232 8192
rect 2296 8128 2304 8192
rect 1904 7104 2304 8128
rect 1904 7040 1912 7104
rect 1976 7040 1992 7104
rect 2056 7040 2072 7104
rect 2136 7040 2152 7104
rect 2216 7040 2232 7104
rect 2296 7040 2304 7104
rect 1904 6016 2304 7040
rect 1904 5952 1912 6016
rect 1976 5952 1992 6016
rect 2056 5952 2072 6016
rect 2136 5952 2152 6016
rect 2216 5952 2232 6016
rect 2296 5952 2304 6016
rect 1904 4928 2304 5952
rect 1904 4864 1912 4928
rect 1976 4864 1992 4928
rect 2056 4864 2072 4928
rect 2136 4864 2152 4928
rect 2216 4864 2232 4928
rect 2296 4864 2304 4928
rect 1904 3840 2304 4864
rect 1904 3776 1912 3840
rect 1976 3776 1992 3840
rect 2056 3776 2072 3840
rect 2136 3776 2152 3840
rect 2216 3776 2232 3840
rect 2296 3776 2304 3840
rect 1904 3294 2304 3776
rect 1904 3058 1986 3294
rect 2222 3058 2304 3294
rect 1904 2752 2304 3058
rect 1904 2688 1912 2752
rect 1976 2688 1992 2752
rect 2056 2688 2072 2752
rect 2136 2688 2152 2752
rect 2216 2688 2232 2752
rect 2296 2688 2304 2752
rect 1904 2128 2304 2688
rect 2644 18528 3044 18544
rect 2644 18464 2652 18528
rect 2716 18464 2732 18528
rect 2796 18464 2812 18528
rect 2876 18464 2892 18528
rect 2956 18464 2972 18528
rect 3036 18464 3044 18528
rect 2644 17440 3044 18464
rect 2644 17376 2652 17440
rect 2716 17376 2732 17440
rect 2796 17376 2812 17440
rect 2876 17376 2892 17440
rect 2956 17376 2972 17440
rect 3036 17376 3044 17440
rect 2644 16352 3044 17376
rect 2644 16288 2652 16352
rect 2716 16288 2732 16352
rect 2796 16288 2812 16352
rect 2876 16288 2892 16352
rect 2956 16288 2972 16352
rect 3036 16288 3044 16352
rect 2644 16034 3044 16288
rect 2644 15798 2726 16034
rect 2962 15798 3044 16034
rect 2644 15264 3044 15798
rect 2644 15200 2652 15264
rect 2716 15200 2732 15264
rect 2796 15200 2812 15264
rect 2876 15200 2892 15264
rect 2956 15200 2972 15264
rect 3036 15200 3044 15264
rect 2644 14176 3044 15200
rect 2644 14112 2652 14176
rect 2716 14112 2732 14176
rect 2796 14112 2812 14176
rect 2876 14112 2892 14176
rect 2956 14112 2972 14176
rect 3036 14112 3044 14176
rect 2644 13088 3044 14112
rect 2644 13024 2652 13088
rect 2716 13024 2732 13088
rect 2796 13024 2812 13088
rect 2876 13024 2892 13088
rect 2956 13024 2972 13088
rect 3036 13024 3044 13088
rect 2644 12000 3044 13024
rect 2644 11936 2652 12000
rect 2716 11936 2732 12000
rect 2796 11936 2812 12000
rect 2876 11936 2892 12000
rect 2956 11936 2972 12000
rect 3036 11936 3044 12000
rect 2644 10912 3044 11936
rect 2644 10848 2652 10912
rect 2716 10848 2732 10912
rect 2796 10848 2812 10912
rect 2876 10848 2892 10912
rect 2956 10848 2972 10912
rect 3036 10848 3044 10912
rect 2644 10034 3044 10848
rect 2644 9824 2726 10034
rect 2962 9824 3044 10034
rect 2644 9760 2652 9824
rect 2716 9798 2726 9824
rect 2962 9798 2972 9824
rect 2716 9760 2732 9798
rect 2796 9760 2812 9798
rect 2876 9760 2892 9798
rect 2956 9760 2972 9798
rect 3036 9760 3044 9824
rect 2644 8736 3044 9760
rect 2644 8672 2652 8736
rect 2716 8672 2732 8736
rect 2796 8672 2812 8736
rect 2876 8672 2892 8736
rect 2956 8672 2972 8736
rect 3036 8672 3044 8736
rect 2644 7648 3044 8672
rect 2644 7584 2652 7648
rect 2716 7584 2732 7648
rect 2796 7584 2812 7648
rect 2876 7584 2892 7648
rect 2956 7584 2972 7648
rect 3036 7584 3044 7648
rect 2644 6560 3044 7584
rect 2644 6496 2652 6560
rect 2716 6496 2732 6560
rect 2796 6496 2812 6560
rect 2876 6496 2892 6560
rect 2956 6496 2972 6560
rect 3036 6496 3044 6560
rect 2644 5472 3044 6496
rect 2644 5408 2652 5472
rect 2716 5408 2732 5472
rect 2796 5408 2812 5472
rect 2876 5408 2892 5472
rect 2956 5408 2972 5472
rect 3036 5408 3044 5472
rect 2644 4384 3044 5408
rect 2644 4320 2652 4384
rect 2716 4320 2732 4384
rect 2796 4320 2812 4384
rect 2876 4320 2892 4384
rect 2956 4320 2972 4384
rect 3036 4320 3044 4384
rect 2644 4034 3044 4320
rect 2644 3798 2726 4034
rect 2962 3798 3044 4034
rect 2644 3296 3044 3798
rect 2644 3232 2652 3296
rect 2716 3232 2732 3296
rect 2796 3232 2812 3296
rect 2876 3232 2892 3296
rect 2956 3232 2972 3296
rect 3036 3232 3044 3296
rect 2644 2208 3044 3232
rect 2644 2144 2652 2208
rect 2716 2144 2732 2208
rect 2796 2144 2812 2208
rect 2876 2144 2892 2208
rect 2956 2144 2972 2208
rect 3036 2144 3044 2208
rect 2644 2128 3044 2144
rect 7904 17984 8304 18544
rect 7904 17920 7912 17984
rect 7976 17920 7992 17984
rect 8056 17920 8072 17984
rect 8136 17920 8152 17984
rect 8216 17920 8232 17984
rect 8296 17920 8304 17984
rect 7904 16896 8304 17920
rect 7904 16832 7912 16896
rect 7976 16832 7992 16896
rect 8056 16832 8072 16896
rect 8136 16832 8152 16896
rect 8216 16832 8232 16896
rect 8296 16832 8304 16896
rect 7904 15808 8304 16832
rect 7904 15744 7912 15808
rect 7976 15744 7992 15808
rect 8056 15744 8072 15808
rect 8136 15744 8152 15808
rect 8216 15744 8232 15808
rect 8296 15744 8304 15808
rect 7904 15294 8304 15744
rect 7904 15058 7986 15294
rect 8222 15058 8304 15294
rect 7904 14720 8304 15058
rect 7904 14656 7912 14720
rect 7976 14656 7992 14720
rect 8056 14656 8072 14720
rect 8136 14656 8152 14720
rect 8216 14656 8232 14720
rect 8296 14656 8304 14720
rect 7904 13632 8304 14656
rect 7904 13568 7912 13632
rect 7976 13568 7992 13632
rect 8056 13568 8072 13632
rect 8136 13568 8152 13632
rect 8216 13568 8232 13632
rect 8296 13568 8304 13632
rect 7904 12544 8304 13568
rect 7904 12480 7912 12544
rect 7976 12480 7992 12544
rect 8056 12480 8072 12544
rect 8136 12480 8152 12544
rect 8216 12480 8232 12544
rect 8296 12480 8304 12544
rect 7904 11456 8304 12480
rect 7904 11392 7912 11456
rect 7976 11392 7992 11456
rect 8056 11392 8072 11456
rect 8136 11392 8152 11456
rect 8216 11392 8232 11456
rect 8296 11392 8304 11456
rect 7904 10368 8304 11392
rect 7904 10304 7912 10368
rect 7976 10304 7992 10368
rect 8056 10304 8072 10368
rect 8136 10304 8152 10368
rect 8216 10304 8232 10368
rect 8296 10304 8304 10368
rect 7904 9294 8304 10304
rect 7904 9280 7986 9294
rect 8222 9280 8304 9294
rect 7904 9216 7912 9280
rect 7976 9216 7986 9280
rect 8222 9216 8232 9280
rect 8296 9216 8304 9280
rect 7904 9058 7986 9216
rect 8222 9058 8304 9216
rect 7904 8192 8304 9058
rect 7904 8128 7912 8192
rect 7976 8128 7992 8192
rect 8056 8128 8072 8192
rect 8136 8128 8152 8192
rect 8216 8128 8232 8192
rect 8296 8128 8304 8192
rect 7904 7104 8304 8128
rect 7904 7040 7912 7104
rect 7976 7040 7992 7104
rect 8056 7040 8072 7104
rect 8136 7040 8152 7104
rect 8216 7040 8232 7104
rect 8296 7040 8304 7104
rect 7904 6016 8304 7040
rect 7904 5952 7912 6016
rect 7976 5952 7992 6016
rect 8056 5952 8072 6016
rect 8136 5952 8152 6016
rect 8216 5952 8232 6016
rect 8296 5952 8304 6016
rect 7904 4928 8304 5952
rect 7904 4864 7912 4928
rect 7976 4864 7992 4928
rect 8056 4864 8072 4928
rect 8136 4864 8152 4928
rect 8216 4864 8232 4928
rect 8296 4864 8304 4928
rect 7904 3840 8304 4864
rect 7904 3776 7912 3840
rect 7976 3776 7992 3840
rect 8056 3776 8072 3840
rect 8136 3776 8152 3840
rect 8216 3776 8232 3840
rect 8296 3776 8304 3840
rect 7904 3294 8304 3776
rect 7904 3058 7986 3294
rect 8222 3058 8304 3294
rect 7904 2752 8304 3058
rect 7904 2688 7912 2752
rect 7976 2688 7992 2752
rect 8056 2688 8072 2752
rect 8136 2688 8152 2752
rect 8216 2688 8232 2752
rect 8296 2688 8304 2752
rect 7904 2128 8304 2688
rect 8644 18528 9044 18544
rect 8644 18464 8652 18528
rect 8716 18464 8732 18528
rect 8796 18464 8812 18528
rect 8876 18464 8892 18528
rect 8956 18464 8972 18528
rect 9036 18464 9044 18528
rect 8644 17440 9044 18464
rect 12571 18052 12637 18053
rect 12571 17988 12572 18052
rect 12636 17988 12637 18052
rect 12571 17987 12637 17988
rect 8644 17376 8652 17440
rect 8716 17376 8732 17440
rect 8796 17376 8812 17440
rect 8876 17376 8892 17440
rect 8956 17376 8972 17440
rect 9036 17376 9044 17440
rect 8644 16352 9044 17376
rect 8644 16288 8652 16352
rect 8716 16288 8732 16352
rect 8796 16288 8812 16352
rect 8876 16288 8892 16352
rect 8956 16288 8972 16352
rect 9036 16288 9044 16352
rect 8644 16034 9044 16288
rect 8644 15798 8726 16034
rect 8962 15798 9044 16034
rect 8644 15264 9044 15798
rect 8644 15200 8652 15264
rect 8716 15200 8732 15264
rect 8796 15200 8812 15264
rect 8876 15200 8892 15264
rect 8956 15200 8972 15264
rect 9036 15200 9044 15264
rect 8644 14176 9044 15200
rect 8644 14112 8652 14176
rect 8716 14112 8732 14176
rect 8796 14112 8812 14176
rect 8876 14112 8892 14176
rect 8956 14112 8972 14176
rect 9036 14112 9044 14176
rect 8644 13088 9044 14112
rect 8644 13024 8652 13088
rect 8716 13024 8732 13088
rect 8796 13024 8812 13088
rect 8876 13024 8892 13088
rect 8956 13024 8972 13088
rect 9036 13024 9044 13088
rect 8644 12000 9044 13024
rect 8644 11936 8652 12000
rect 8716 11936 8732 12000
rect 8796 11936 8812 12000
rect 8876 11936 8892 12000
rect 8956 11936 8972 12000
rect 9036 11936 9044 12000
rect 8644 10912 9044 11936
rect 8644 10848 8652 10912
rect 8716 10848 8732 10912
rect 8796 10848 8812 10912
rect 8876 10848 8892 10912
rect 8956 10848 8972 10912
rect 9036 10848 9044 10912
rect 8644 10034 9044 10848
rect 8644 9824 8726 10034
rect 8962 9824 9044 10034
rect 8644 9760 8652 9824
rect 8716 9798 8726 9824
rect 8962 9798 8972 9824
rect 8716 9760 8732 9798
rect 8796 9760 8812 9798
rect 8876 9760 8892 9798
rect 8956 9760 8972 9798
rect 9036 9760 9044 9824
rect 8644 8736 9044 9760
rect 8644 8672 8652 8736
rect 8716 8672 8732 8736
rect 8796 8672 8812 8736
rect 8876 8672 8892 8736
rect 8956 8672 8972 8736
rect 9036 8672 9044 8736
rect 8644 7648 9044 8672
rect 12574 7717 12634 17987
rect 13904 17984 14304 18544
rect 13904 17920 13912 17984
rect 13976 17920 13992 17984
rect 14056 17920 14072 17984
rect 14136 17920 14152 17984
rect 14216 17920 14232 17984
rect 14296 17920 14304 17984
rect 13904 16896 14304 17920
rect 13904 16832 13912 16896
rect 13976 16832 13992 16896
rect 14056 16832 14072 16896
rect 14136 16832 14152 16896
rect 14216 16832 14232 16896
rect 14296 16832 14304 16896
rect 13904 15808 14304 16832
rect 13904 15744 13912 15808
rect 13976 15744 13992 15808
rect 14056 15744 14072 15808
rect 14136 15744 14152 15808
rect 14216 15744 14232 15808
rect 14296 15744 14304 15808
rect 13904 15294 14304 15744
rect 13904 15058 13986 15294
rect 14222 15058 14304 15294
rect 13904 14720 14304 15058
rect 13904 14656 13912 14720
rect 13976 14656 13992 14720
rect 14056 14656 14072 14720
rect 14136 14656 14152 14720
rect 14216 14656 14232 14720
rect 14296 14656 14304 14720
rect 13904 13632 14304 14656
rect 13904 13568 13912 13632
rect 13976 13568 13992 13632
rect 14056 13568 14072 13632
rect 14136 13568 14152 13632
rect 14216 13568 14232 13632
rect 14296 13568 14304 13632
rect 13904 12544 14304 13568
rect 13904 12480 13912 12544
rect 13976 12480 13992 12544
rect 14056 12480 14072 12544
rect 14136 12480 14152 12544
rect 14216 12480 14232 12544
rect 14296 12480 14304 12544
rect 13904 11456 14304 12480
rect 13904 11392 13912 11456
rect 13976 11392 13992 11456
rect 14056 11392 14072 11456
rect 14136 11392 14152 11456
rect 14216 11392 14232 11456
rect 14296 11392 14304 11456
rect 13904 10368 14304 11392
rect 13904 10304 13912 10368
rect 13976 10304 13992 10368
rect 14056 10304 14072 10368
rect 14136 10304 14152 10368
rect 14216 10304 14232 10368
rect 14296 10304 14304 10368
rect 13904 9294 14304 10304
rect 14644 18528 15044 18544
rect 14644 18464 14652 18528
rect 14716 18464 14732 18528
rect 14796 18464 14812 18528
rect 14876 18464 14892 18528
rect 14956 18464 14972 18528
rect 15036 18464 15044 18528
rect 14644 17440 15044 18464
rect 14644 17376 14652 17440
rect 14716 17376 14732 17440
rect 14796 17376 14812 17440
rect 14876 17376 14892 17440
rect 14956 17376 14972 17440
rect 15036 17376 15044 17440
rect 14644 16352 15044 17376
rect 14644 16288 14652 16352
rect 14716 16288 14732 16352
rect 14796 16288 14812 16352
rect 14876 16288 14892 16352
rect 14956 16288 14972 16352
rect 15036 16288 15044 16352
rect 14644 16034 15044 16288
rect 14644 15798 14726 16034
rect 14962 15798 15044 16034
rect 14644 15264 15044 15798
rect 14644 15200 14652 15264
rect 14716 15200 14732 15264
rect 14796 15200 14812 15264
rect 14876 15200 14892 15264
rect 14956 15200 14972 15264
rect 15036 15200 15044 15264
rect 14644 14176 15044 15200
rect 14644 14112 14652 14176
rect 14716 14112 14732 14176
rect 14796 14112 14812 14176
rect 14876 14112 14892 14176
rect 14956 14112 14972 14176
rect 15036 14112 15044 14176
rect 14644 13088 15044 14112
rect 14644 13024 14652 13088
rect 14716 13024 14732 13088
rect 14796 13024 14812 13088
rect 14876 13024 14892 13088
rect 14956 13024 14972 13088
rect 15036 13024 15044 13088
rect 14644 12000 15044 13024
rect 14644 11936 14652 12000
rect 14716 11936 14732 12000
rect 14796 11936 14812 12000
rect 14876 11936 14892 12000
rect 14956 11936 14972 12000
rect 15036 11936 15044 12000
rect 14644 10912 15044 11936
rect 14644 10848 14652 10912
rect 14716 10848 14732 10912
rect 14796 10848 14812 10912
rect 14876 10848 14892 10912
rect 14956 10848 14972 10912
rect 15036 10848 15044 10912
rect 14644 10034 15044 10848
rect 14644 9824 14726 10034
rect 14962 9824 15044 10034
rect 14644 9760 14652 9824
rect 14716 9798 14726 9824
rect 14962 9798 14972 9824
rect 14716 9760 14732 9798
rect 14796 9760 14812 9798
rect 14876 9760 14892 9798
rect 14956 9760 14972 9798
rect 15036 9760 15044 9824
rect 14411 9484 14477 9485
rect 14411 9420 14412 9484
rect 14476 9420 14477 9484
rect 14411 9419 14477 9420
rect 13904 9280 13986 9294
rect 14222 9280 14304 9294
rect 13904 9216 13912 9280
rect 13976 9216 13986 9280
rect 14222 9216 14232 9280
rect 14296 9216 14304 9280
rect 13904 9058 13986 9216
rect 14222 9058 14304 9216
rect 13904 8192 14304 9058
rect 13904 8128 13912 8192
rect 13976 8128 13992 8192
rect 14056 8128 14072 8192
rect 14136 8128 14152 8192
rect 14216 8128 14232 8192
rect 14296 8128 14304 8192
rect 12571 7716 12637 7717
rect 12571 7652 12572 7716
rect 12636 7652 12637 7716
rect 12571 7651 12637 7652
rect 8644 7584 8652 7648
rect 8716 7584 8732 7648
rect 8796 7584 8812 7648
rect 8876 7584 8892 7648
rect 8956 7584 8972 7648
rect 9036 7584 9044 7648
rect 8644 6560 9044 7584
rect 8644 6496 8652 6560
rect 8716 6496 8732 6560
rect 8796 6496 8812 6560
rect 8876 6496 8892 6560
rect 8956 6496 8972 6560
rect 9036 6496 9044 6560
rect 8644 5472 9044 6496
rect 8644 5408 8652 5472
rect 8716 5408 8732 5472
rect 8796 5408 8812 5472
rect 8876 5408 8892 5472
rect 8956 5408 8972 5472
rect 9036 5408 9044 5472
rect 8644 4384 9044 5408
rect 8644 4320 8652 4384
rect 8716 4320 8732 4384
rect 8796 4320 8812 4384
rect 8876 4320 8892 4384
rect 8956 4320 8972 4384
rect 9036 4320 9044 4384
rect 8644 4034 9044 4320
rect 8644 3798 8726 4034
rect 8962 3798 9044 4034
rect 8644 3296 9044 3798
rect 8644 3232 8652 3296
rect 8716 3232 8732 3296
rect 8796 3232 8812 3296
rect 8876 3232 8892 3296
rect 8956 3232 8972 3296
rect 9036 3232 9044 3296
rect 8644 2208 9044 3232
rect 8644 2144 8652 2208
rect 8716 2144 8732 2208
rect 8796 2144 8812 2208
rect 8876 2144 8892 2208
rect 8956 2144 8972 2208
rect 9036 2144 9044 2208
rect 8644 2128 9044 2144
rect 13904 7104 14304 8128
rect 13904 7040 13912 7104
rect 13976 7040 13992 7104
rect 14056 7040 14072 7104
rect 14136 7040 14152 7104
rect 14216 7040 14232 7104
rect 14296 7040 14304 7104
rect 13904 6016 14304 7040
rect 14414 6493 14474 9419
rect 14644 8736 15044 9760
rect 14644 8672 14652 8736
rect 14716 8672 14732 8736
rect 14796 8672 14812 8736
rect 14876 8672 14892 8736
rect 14956 8672 14972 8736
rect 15036 8672 15044 8736
rect 14644 7648 15044 8672
rect 14644 7584 14652 7648
rect 14716 7584 14732 7648
rect 14796 7584 14812 7648
rect 14876 7584 14892 7648
rect 14956 7584 14972 7648
rect 15036 7584 15044 7648
rect 14644 6560 15044 7584
rect 14644 6496 14652 6560
rect 14716 6496 14732 6560
rect 14796 6496 14812 6560
rect 14876 6496 14892 6560
rect 14956 6496 14972 6560
rect 15036 6496 15044 6560
rect 14411 6492 14477 6493
rect 14411 6428 14412 6492
rect 14476 6428 14477 6492
rect 14411 6427 14477 6428
rect 13904 5952 13912 6016
rect 13976 5952 13992 6016
rect 14056 5952 14072 6016
rect 14136 5952 14152 6016
rect 14216 5952 14232 6016
rect 14296 5952 14304 6016
rect 13904 4928 14304 5952
rect 13904 4864 13912 4928
rect 13976 4864 13992 4928
rect 14056 4864 14072 4928
rect 14136 4864 14152 4928
rect 14216 4864 14232 4928
rect 14296 4864 14304 4928
rect 13904 3840 14304 4864
rect 13904 3776 13912 3840
rect 13976 3776 13992 3840
rect 14056 3776 14072 3840
rect 14136 3776 14152 3840
rect 14216 3776 14232 3840
rect 14296 3776 14304 3840
rect 13904 3294 14304 3776
rect 13904 3058 13986 3294
rect 14222 3058 14304 3294
rect 13904 2752 14304 3058
rect 13904 2688 13912 2752
rect 13976 2688 13992 2752
rect 14056 2688 14072 2752
rect 14136 2688 14152 2752
rect 14216 2688 14232 2752
rect 14296 2688 14304 2752
rect 13904 2128 14304 2688
rect 14644 5472 15044 6496
rect 14644 5408 14652 5472
rect 14716 5408 14732 5472
rect 14796 5408 14812 5472
rect 14876 5408 14892 5472
rect 14956 5408 14972 5472
rect 15036 5408 15044 5472
rect 14644 4384 15044 5408
rect 14644 4320 14652 4384
rect 14716 4320 14732 4384
rect 14796 4320 14812 4384
rect 14876 4320 14892 4384
rect 14956 4320 14972 4384
rect 15036 4320 15044 4384
rect 14644 4034 15044 4320
rect 14644 3798 14726 4034
rect 14962 3798 15044 4034
rect 14644 3296 15044 3798
rect 14644 3232 14652 3296
rect 14716 3232 14732 3296
rect 14796 3232 14812 3296
rect 14876 3232 14892 3296
rect 14956 3232 14972 3296
rect 15036 3232 15044 3296
rect 14644 2208 15044 3232
rect 14644 2144 14652 2208
rect 14716 2144 14732 2208
rect 14796 2144 14812 2208
rect 14876 2144 14892 2208
rect 14956 2144 14972 2208
rect 15036 2144 15044 2208
rect 14644 2128 15044 2144
<< via4 >>
rect 1986 15058 2222 15294
rect 1986 9280 2222 9294
rect 1986 9216 1992 9280
rect 1992 9216 2056 9280
rect 2056 9216 2072 9280
rect 2072 9216 2136 9280
rect 2136 9216 2152 9280
rect 2152 9216 2216 9280
rect 2216 9216 2222 9280
rect 1986 9058 2222 9216
rect 1986 3058 2222 3294
rect 2726 15798 2962 16034
rect 2726 9824 2962 10034
rect 2726 9798 2732 9824
rect 2732 9798 2796 9824
rect 2796 9798 2812 9824
rect 2812 9798 2876 9824
rect 2876 9798 2892 9824
rect 2892 9798 2956 9824
rect 2956 9798 2962 9824
rect 2726 3798 2962 4034
rect 7986 15058 8222 15294
rect 7986 9280 8222 9294
rect 7986 9216 7992 9280
rect 7992 9216 8056 9280
rect 8056 9216 8072 9280
rect 8072 9216 8136 9280
rect 8136 9216 8152 9280
rect 8152 9216 8216 9280
rect 8216 9216 8222 9280
rect 7986 9058 8222 9216
rect 7986 3058 8222 3294
rect 8726 15798 8962 16034
rect 8726 9824 8962 10034
rect 8726 9798 8732 9824
rect 8732 9798 8796 9824
rect 8796 9798 8812 9824
rect 8812 9798 8876 9824
rect 8876 9798 8892 9824
rect 8892 9798 8956 9824
rect 8956 9798 8962 9824
rect 13986 15058 14222 15294
rect 14726 15798 14962 16034
rect 14726 9824 14962 10034
rect 14726 9798 14732 9824
rect 14732 9798 14796 9824
rect 14796 9798 14812 9824
rect 14812 9798 14876 9824
rect 14876 9798 14892 9824
rect 14892 9798 14956 9824
rect 14956 9798 14962 9824
rect 13986 9280 14222 9294
rect 13986 9216 13992 9280
rect 13992 9216 14056 9280
rect 14056 9216 14072 9280
rect 14072 9216 14136 9280
rect 14136 9216 14152 9280
rect 14152 9216 14216 9280
rect 14216 9216 14222 9280
rect 13986 9058 14222 9216
rect 8726 3798 8962 4034
rect 13986 3058 14222 3294
rect 14726 3798 14962 4034
<< metal5 >>
rect 1056 16034 17896 16116
rect 1056 15798 2726 16034
rect 2962 15798 8726 16034
rect 8962 15798 14726 16034
rect 14962 15798 17896 16034
rect 1056 15716 17896 15798
rect 1056 15294 17896 15376
rect 1056 15058 1986 15294
rect 2222 15058 7986 15294
rect 8222 15058 13986 15294
rect 14222 15058 17896 15294
rect 1056 14976 17896 15058
rect 1056 10034 17896 10116
rect 1056 9798 2726 10034
rect 2962 9798 8726 10034
rect 8962 9798 14726 10034
rect 14962 9798 17896 10034
rect 1056 9716 17896 9798
rect 1056 9294 17896 9376
rect 1056 9058 1986 9294
rect 2222 9058 7986 9294
rect 8222 9058 13986 9294
rect 14222 9058 17896 9294
rect 1056 8976 17896 9058
rect 1056 4034 17896 4116
rect 1056 3798 2726 4034
rect 2962 3798 8726 4034
rect 8962 3798 14726 4034
rect 14962 3798 17896 4034
rect 1056 3716 17896 3798
rect 1056 3294 17896 3376
rect 1056 3058 1986 3294
rect 2222 3058 7986 3294
rect 8222 3058 13986 3294
rect 14222 3058 17896 3294
rect 1056 2976 17896 3058
use sky130_fd_sc_hd__inv_2  _313_
timestamp 1
transform 1 0 17112 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _314_
timestamp 1
transform 1 0 14260 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _315_
timestamp 1
transform 1 0 13340 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _316_
timestamp 1
transform 1 0 14168 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _317_
timestamp 1
transform 1 0 13064 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _318_
timestamp 1
transform -1 0 4048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _319_
timestamp 1
transform -1 0 3496 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _320_
timestamp 1
transform -1 0 7728 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _321_
timestamp 1
transform 1 0 7360 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _322_
timestamp 1
transform -1 0 7360 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _323_
timestamp 1
transform 1 0 11868 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _324_
timestamp 1
transform 1 0 8556 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _325_
timestamp 1
transform 1 0 7268 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _326_
timestamp 1
transform 1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _327_
timestamp 1
transform 1 0 7452 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _328_
timestamp 1
transform -1 0 8188 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _329_
timestamp 1
transform 1 0 7912 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _330_
timestamp 1
transform -1 0 8740 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _331_
timestamp 1
transform 1 0 13064 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_4  _332_
timestamp 1
transform 1 0 13064 0 -1 3264
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _333_
timestamp 1
transform -1 0 11224 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _334_
timestamp 1
transform 1 0 8832 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _335_
timestamp 1
transform -1 0 8832 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _336_
timestamp 1
transform -1 0 8280 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _337_
timestamp 1
transform -1 0 10580 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _338_
timestamp 1
transform -1 0 10028 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor3b_1  _339_
timestamp 1
transform 1 0 13432 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _340_
timestamp 1
transform -1 0 13064 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _341_
timestamp 1
transform 1 0 8924 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _342_
timestamp 1
transform 1 0 7728 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _343_
timestamp 1
transform 1 0 6992 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _344_
timestamp 1
transform 1 0 12696 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _345_
timestamp 1
transform 1 0 12236 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _346_
timestamp 1
transform 1 0 11500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _347_
timestamp 1
transform 1 0 15640 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _348_
timestamp 1
transform 1 0 12972 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _349_
timestamp 1
transform 1 0 12052 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _350_
timestamp 1
transform -1 0 6440 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _351_
timestamp 1
transform 1 0 6992 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _352_
timestamp 1
transform -1 0 6992 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _353_
timestamp 1
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _354_
timestamp 1
transform -1 0 6532 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _355_
timestamp 1
transform -1 0 4876 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _356_
timestamp 1
transform -1 0 4324 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _357_
timestamp 1
transform -1 0 17112 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _358_
timestamp 1
transform -1 0 16560 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _359_
timestamp 1
transform -1 0 17388 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _360_
timestamp 1
transform 1 0 16376 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _361_
timestamp 1
transform 1 0 16652 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_2  _362_
timestamp 1
transform 1 0 16192 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _363_
timestamp 1
transform 1 0 17020 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _364_
timestamp 1
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _365_
timestamp 1
transform 1 0 16652 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _366_
timestamp 1
transform 1 0 8188 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _367_
timestamp 1
transform 1 0 8924 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _368_
timestamp 1
transform 1 0 10672 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _369_
timestamp 1
transform -1 0 11316 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o221ai_2  _370_
timestamp 1
transform 1 0 10580 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__or3_1  _371_
timestamp 1
transform -1 0 11316 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_1  _372_
timestamp 1
transform 1 0 10488 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _373_
timestamp 1
transform 1 0 10120 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _374_
timestamp 1
transform -1 0 9568 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _375_
timestamp 1
transform -1 0 10764 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _376_
timestamp 1
transform -1 0 10488 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _377_
timestamp 1
transform 1 0 9844 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _378_
timestamp 1
transform -1 0 5980 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _379_
timestamp 1
transform 1 0 4968 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _380_
timestamp 1
transform -1 0 4784 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _381_
timestamp 1
transform -1 0 4140 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _382_
timestamp 1
transform -1 0 16560 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_2  _383_
timestamp 1
transform 1 0 16652 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _384_
timestamp 1
transform 1 0 16192 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _385_
timestamp 1
transform 1 0 16100 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _386_
timestamp 1
transform -1 0 15364 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _387_
timestamp 1
transform 1 0 16652 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _388_
timestamp 1
transform -1 0 17112 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _389_
timestamp 1
transform -1 0 15548 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _390_
timestamp 1
transform -1 0 12420 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _391_
timestamp 1
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _392_
timestamp 1
transform -1 0 15732 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _393_
timestamp 1
transform 1 0 15088 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _394_
timestamp 1
transform -1 0 15640 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _395_
timestamp 1
transform -1 0 17296 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _396_
timestamp 1
transform 1 0 16008 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _397_
timestamp 1
transform 1 0 16100 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _398_
timestamp 1
transform 1 0 15732 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _399_
timestamp 1
transform -1 0 17020 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _400_
timestamp 1
transform -1 0 10304 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _401_
timestamp 1
transform -1 0 6256 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _402_
timestamp 1
transform -1 0 6992 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _403_
timestamp 1
transform -1 0 6716 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _404_
timestamp 1
transform -1 0 6164 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _405_
timestamp 1
transform 1 0 4232 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _406_
timestamp 1
transform -1 0 4232 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _407_
timestamp 1
transform -1 0 15640 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _408_
timestamp 1
transform -1 0 15916 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _409_
timestamp 1
transform -1 0 15180 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _410_
timestamp 1
transform 1 0 15640 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _411_
timestamp 1
transform 1 0 14904 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _412_
timestamp 1
transform -1 0 15640 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _413_
timestamp 1
transform -1 0 15088 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _414_
timestamp 1
transform -1 0 9200 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _415_
timestamp 1
transform -1 0 13984 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _416_
timestamp 1
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _417_
timestamp 1
transform -1 0 14904 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _418_
timestamp 1
transform 1 0 14628 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _419_
timestamp 1
transform -1 0 15364 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _420_
timestamp 1
transform -1 0 14904 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _421_
timestamp 1
transform 1 0 14352 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _422_
timestamp 1
transform 1 0 14996 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _423_
timestamp 1
transform -1 0 17296 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _424_
timestamp 1
transform 1 0 15732 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _425_
timestamp 1
transform 1 0 16652 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _426_
timestamp 1
transform -1 0 16744 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _427_
timestamp 1
transform -1 0 17572 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _428_
timestamp 1
transform 1 0 4692 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _429_
timestamp 1
transform -1 0 4692 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _430_
timestamp 1
transform -1 0 4784 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _431_
timestamp 1
transform -1 0 4048 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _432_
timestamp 1
transform -1 0 4324 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _433_
timestamp 1
transform -1 0 14904 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _434_
timestamp 1
transform 1 0 14168 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _435_
timestamp 1
transform 1 0 12604 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _436_
timestamp 1
transform -1 0 12696 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _437_
timestamp 1
transform 1 0 15180 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _438_
timestamp 1
transform -1 0 14904 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _439_
timestamp 1
transform 1 0 13708 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _440_
timestamp 1
transform -1 0 15180 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _441_
timestamp 1
transform -1 0 15180 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _442_
timestamp 1
transform -1 0 14444 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _443_
timestamp 1
transform -1 0 12604 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _444_
timestamp 1
transform 1 0 12052 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _445_
timestamp 1
transform 1 0 14352 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _446_
timestamp 1
transform -1 0 9476 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _447_
timestamp 1
transform 1 0 11040 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _448_
timestamp 1
transform -1 0 10304 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _449_
timestamp 1
transform 1 0 13064 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _450_
timestamp 1
transform -1 0 12420 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _451_
timestamp 1
transform 1 0 12420 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _452_
timestamp 1
transform -1 0 10028 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _453_
timestamp 1
transform -1 0 10488 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _454_
timestamp 1
transform 1 0 8924 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _455_
timestamp 1
transform -1 0 15916 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _456_
timestamp 1
transform 1 0 15088 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _457_
timestamp 1
transform 1 0 14536 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _458_
timestamp 1
transform 1 0 14076 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _459_
timestamp 1
transform -1 0 9936 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _460_
timestamp 1
transform -1 0 8280 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _461_
timestamp 1
transform -1 0 7820 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _462_
timestamp 1
transform 1 0 6624 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _463_
timestamp 1
transform 1 0 11684 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _464_
timestamp 1
transform -1 0 7452 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _465_
timestamp 1
transform -1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _466_
timestamp 1
transform 1 0 4968 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _467_
timestamp 1
transform -1 0 5704 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _468_
timestamp 1
transform -1 0 6348 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _469_
timestamp 1
transform -1 0 3496 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _470_
timestamp 1
transform -1 0 13156 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _471_
timestamp 1
transform 1 0 12880 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _472_
timestamp 1
transform -1 0 14076 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _473_
timestamp 1
transform 1 0 15548 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _474_
timestamp 1
transform -1 0 15548 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _475_
timestamp 1
transform 1 0 13340 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_2  _476_
timestamp 1
transform 1 0 11500 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _477_
timestamp 1
transform 1 0 14904 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _478_
timestamp 1
transform 1 0 14444 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _479_
timestamp 1
transform 1 0 14076 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _480_
timestamp 1
transform 1 0 9844 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _481_
timestamp 1
transform -1 0 11960 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _482_
timestamp 1
transform 1 0 9568 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _483_
timestamp 1
transform -1 0 10856 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _484_
timestamp 1
transform 1 0 9200 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _485_
timestamp 1
transform 1 0 7728 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _486_
timestamp 1
transform 1 0 9016 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _487_
timestamp 1
transform -1 0 8740 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _488_
timestamp 1
transform -1 0 9016 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _489_
timestamp 1
transform 1 0 7452 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _490_
timestamp 1
transform 1 0 7084 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _491_
timestamp 1
transform -1 0 7084 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _492_
timestamp 1
transform 1 0 4508 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _493_
timestamp 1
transform -1 0 5520 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _494_
timestamp 1
transform 1 0 4508 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _495_
timestamp 1
transform 1 0 3772 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _496_
timestamp 1
transform -1 0 3864 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _497_
timestamp 1
transform -1 0 4324 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _498_
timestamp 1
transform -1 0 13340 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _499_
timestamp 1
transform -1 0 13064 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _500_
timestamp 1
transform -1 0 13064 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_2  _501_
timestamp 1
transform 1 0 10304 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _502_
timestamp 1
transform 1 0 14076 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _503_
timestamp 1
transform -1 0 12972 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _504_
timestamp 1
transform 1 0 12512 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _505_
timestamp 1
transform 1 0 10212 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _506_
timestamp 1
transform -1 0 14444 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _507_
timestamp 1
transform 1 0 15180 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _508_
timestamp 1
transform 1 0 14444 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _509_
timestamp 1
transform -1 0 11408 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _510_
timestamp 1
transform 1 0 8188 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _511_
timestamp 1
transform 1 0 8556 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _512_
timestamp 1
transform 1 0 8004 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _513_
timestamp 1
transform -1 0 9568 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _514_
timestamp 1
transform 1 0 6900 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _515_
timestamp 1
transform -1 0 7268 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _516_
timestamp 1
transform -1 0 5612 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _517_
timestamp 1
transform -1 0 5336 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _518_
timestamp 1
transform 1 0 4600 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _519_
timestamp 1
transform 1 0 3864 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _520_
timestamp 1
transform 1 0 4324 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _521_
timestamp 1
transform -1 0 4416 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _522_
timestamp 1
transform 1 0 11132 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _523_
timestamp 1
transform -1 0 11592 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _524_
timestamp 1
transform -1 0 15640 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _525_
timestamp 1
transform -1 0 15916 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _526_
timestamp 1
transform 1 0 15824 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _527_
timestamp 1
transform -1 0 15180 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _528_
timestamp 1
transform -1 0 10212 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _529_
timestamp 1
transform 1 0 11040 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _530_
timestamp 1
transform -1 0 11316 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _531_
timestamp 1
transform -1 0 10856 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _532_
timestamp 1
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _533_
timestamp 1
transform 1 0 10120 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _534_
timestamp 1
transform 1 0 7360 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _535_
timestamp 1
transform -1 0 12236 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _536_
timestamp 1
transform 1 0 12236 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _537_
timestamp 1
transform 1 0 13064 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _538_
timestamp 1
transform -1 0 8648 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _539_
timestamp 1
transform -1 0 7636 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _540_
timestamp 1
transform -1 0 7084 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _541_
timestamp 1
transform 1 0 5888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _542_
timestamp 1
transform -1 0 6440 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _543_
timestamp 1
transform -1 0 4968 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _544_
timestamp 1
transform 1 0 3128 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _545_
timestamp 1
transform -1 0 4324 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _546_
timestamp 1
transform 1 0 3312 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _547_
timestamp 1
transform 1 0 3404 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _548_
timestamp 1
transform 1 0 8924 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _549_
timestamp 1
transform -1 0 8556 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _550_
timestamp 1
transform 1 0 13892 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _551_
timestamp 1
transform 1 0 14996 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _552_
timestamp 1
transform -1 0 14996 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a32oi_4  _553_
timestamp 1
transform 1 0 14076 0 1 13056
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _554_
timestamp 1
transform -1 0 9936 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _555_
timestamp 1
transform 1 0 10396 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _556_
timestamp 1
transform 1 0 10396 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _557_
timestamp 1
transform 1 0 11040 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _558_
timestamp 1
transform -1 0 10764 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _559_
timestamp 1
transform 1 0 12788 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _560_
timestamp 1
transform -1 0 12880 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _561_
timestamp 1
transform 1 0 11960 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _562_
timestamp 1
transform -1 0 10396 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _563_
timestamp 1
transform -1 0 6808 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _564_
timestamp 1
transform -1 0 6992 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _565_
timestamp 1
transform 1 0 6348 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _566_
timestamp 1
transform -1 0 6348 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _567_
timestamp 1
transform -1 0 5336 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _568_
timestamp 1
transform -1 0 3496 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _569_
timestamp 1
transform -1 0 15364 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _570_
timestamp 1
transform -1 0 14996 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _571_
timestamp 1
transform -1 0 14168 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _572_
timestamp 1
transform 1 0 12236 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _573_
timestamp 1
transform -1 0 11684 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _574_
timestamp 1
transform -1 0 11408 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _575_
timestamp 1
transform 1 0 9936 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _576_
timestamp 1
transform -1 0 8648 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _577_
timestamp 1
transform -1 0 10488 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _578_
timestamp 1
transform -1 0 7912 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _579_
timestamp 1
transform -1 0 7728 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _580_
timestamp 1
transform -1 0 7176 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _581_
timestamp 1
transform 1 0 5612 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _582_
timestamp 1
transform -1 0 6348 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _583_
timestamp 1
transform -1 0 5612 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _584_
timestamp 1
transform 1 0 4968 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _585_
timestamp 1
transform -1 0 4784 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _586_
timestamp 1
transform -1 0 5704 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _587_
timestamp 1
transform -1 0 4692 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _588_
timestamp 1
transform 1 0 4692 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _589_
timestamp 1
transform 1 0 3956 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _590_
timestamp 1
transform 1 0 12696 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _591_
timestamp 1
transform 1 0 12144 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _592_
timestamp 1
transform 1 0 12972 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _593_
timestamp 1
transform -1 0 8924 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _594_
timestamp 1
transform 1 0 8648 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _595_
timestamp 1
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _596_
timestamp 1
transform 1 0 7820 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _597_
timestamp 1
transform -1 0 6624 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _598_
timestamp 1
transform -1 0 7084 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _599_
timestamp 1
transform -1 0 4876 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _600_
timestamp 1
transform 1 0 4232 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _601_
timestamp 1
transform -1 0 4416 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _602_
timestamp 1
transform 1 0 12880 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _603_
timestamp 1
transform -1 0 7268 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _604_
timestamp 1
transform -1 0 7544 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _605_
timestamp 1
transform -1 0 6808 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _606_
timestamp 1
transform -1 0 6072 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _607_
timestamp 1
transform -1 0 5796 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _608_
timestamp 1
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _609_
timestamp 1
transform 1 0 2852 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _610_
timestamp 1
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _611_
timestamp 1
transform 1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _612_
timestamp 1
transform 1 0 2116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _613_
timestamp 1
transform -1 0 3496 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _614_
timestamp 1
transform -1 0 2484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _615_
timestamp 1
transform -1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _616_
timestamp 1
transform -1 0 2484 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _617_
timestamp 1
transform 1 0 2116 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _618_
timestamp 1
transform -1 0 2576 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _619_
timestamp 1
transform -1 0 3496 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _620_
timestamp 1
transform 1 0 2116 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _621_
timestamp 1
transform -1 0 2484 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _622_
timestamp 1
transform -1 0 2576 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _623_
timestamp 1
transform 1 0 2116 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _624_
timestamp 1
transform -1 0 4048 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _625_
timestamp 1
transform -1 0 4600 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _626_
timestamp 1
transform 1 0 2116 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _627_
timestamp 1
transform 1 0 6532 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _628_
timestamp 1
transform -1 0 6624 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _629_
timestamp 1
transform 1 0 6992 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _630_
timestamp 1
transform -1 0 9200 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _631_
timestamp 1
transform 1 0 12420 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _632_
timestamp 1
transform -1 0 9292 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _633_
timestamp 1
transform 1 0 10856 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _634_
timestamp 1
transform -1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _635_
timestamp 1
transform -1 0 12604 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _636_
timestamp 1
transform -1 0 13524 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _637_
timestamp 1
transform -1 0 14352 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _638_
timestamp 1
transform 1 0 16652 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _639_
timestamp 1
transform 1 0 15548 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _640_
timestamp 1
transform 1 0 16836 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _641_
timestamp 1
transform 1 0 16836 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _642_
timestamp 1
transform -1 0 4232 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _643_
timestamp 1
transform -1 0 6072 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _644_
timestamp 1
transform -1 0 3220 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _645_
timestamp 1
transform -1 0 3220 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _646_
timestamp 1
transform -1 0 3220 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _647_
timestamp 1
transform -1 0 3220 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _648_
timestamp 1
transform -1 0 3220 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _649_
timestamp 1
transform -1 0 3220 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _650_
timestamp 1
transform -1 0 3220 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _651_
timestamp 1
transform -1 0 3220 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _652_
timestamp 1
transform -1 0 3220 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _653_
timestamp 1
transform -1 0 3220 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _654_
timestamp 1
transform -1 0 3220 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _655_
timestamp 1
transform -1 0 3220 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _656_
timestamp 1
transform -1 0 4692 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _657_
timestamp 1
transform -1 0 5336 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _658_
timestamp 1
transform 1 0 1380 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _659_
timestamp 1
transform 1 0 6348 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _660_
timestamp 1
transform 1 0 4600 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _661_
timestamp 1
transform 1 0 6348 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _662_
timestamp 1
transform 1 0 6716 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _663_
timestamp 1
transform 1 0 11868 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _664_
timestamp 1
transform 1 0 7912 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _665_
timestamp 1
transform 1 0 9844 0 1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _666_
timestamp 1
transform 1 0 9752 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _667_
timestamp 1
transform 1 0 11040 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _668_
timestamp 1
transform 1 0 12144 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _669_
timestamp 1
transform 1 0 12972 0 -1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _670_
timestamp 1
transform 1 0 15640 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _671_
timestamp 1
transform 1 0 14628 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _672_
timestamp 1
transform 1 0 15732 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _673_
timestamp 1
transform -1 0 17572 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1
transform -1 0 11316 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1
transform -1 0 8188 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1
transform -1 0 8188 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1
transform 1 0 8832 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1
transform 1 0 11960 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  clkload0
timestamp 1
transform 1 0 5704 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__bufinv_16  clkload1
timestamp 1
transform 1 0 8924 0 1 13056
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_2  clkload2
timestamp 1
transform -1 0 11960 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23
timestamp 1
transform 1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 1
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32
timestamp 1636968456
transform 1 0 4048 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44
timestamp 1
transform 1 0 5152 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48
timestamp 1
transform 1 0 5520 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636968456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636968456
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85
timestamp 1
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636968456
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125
timestamp 1
transform 1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_129
timestamp 1
transform 1 0 12972 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_133
timestamp 1
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636968456
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636968456
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_177
timestamp 1
transform 1 0 17388 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_6
timestamp 1
transform 1 0 1656 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_10
timestamp 1
transform 1 0 2024 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_71
timestamp 1
transform 1 0 7636 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_1_90
timestamp 1
transform 1 0 9384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_119
timestamp 1
transform 1 0 12052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_159
timestamp 1
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_169
timestamp 1
transform 1 0 16652 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_177
timestamp 1
transform 1 0 17388 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_6
timestamp 1636968456
transform 1 0 1656 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_18
timestamp 1
transform 1 0 2760 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636968456
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_41
timestamp 1
transform 1 0 4876 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_49
timestamp 1
transform 1 0 5612 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_59
timestamp 1
transform 1 0 6532 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_67
timestamp 1
transform 1 0 7268 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_72
timestamp 1
transform 1 0 7728 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_92
timestamp 1
transform 1 0 9568 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_100
timestamp 1
transform 1 0 10304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_115
timestamp 1
transform 1 0 11684 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_135
timestamp 1
transform 1 0 13524 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_163
timestamp 1636968456
transform 1 0 16100 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_175
timestamp 1
transform 1 0 17204 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_26
timestamp 1
transform 1 0 3496 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_41
timestamp 1
transform 1 0 4876 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_49
timestamp 1
transform 1 0 5612 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_67
timestamp 1
transform 1 0 7268 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_75
timestamp 1
transform 1 0 8004 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_83
timestamp 1636968456
transform 1 0 8740 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_95
timestamp 1
transform 1 0 9844 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_103
timestamp 1
transform 1 0 10580 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_113
timestamp 1
transform 1 0 11500 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_140
timestamp 1
transform 1 0 13984 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_146
timestamp 1
transform 1 0 14536 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_159
timestamp 1
transform 1 0 15732 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_169
timestamp 1
transform 1 0 16652 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_177
timestamp 1
transform 1 0 17388 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_6
timestamp 1
transform 1 0 1656 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636968456
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636968456
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636968456
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_53
timestamp 1
transform 1 0 5980 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_58
timestamp 1636968456
transform 1 0 6440 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_70
timestamp 1636968456
transform 1 0 7544 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_94
timestamp 1
transform 1 0 9752 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_111
timestamp 1636968456
transform 1 0 11316 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_123
timestamp 1636968456
transform 1 0 12420 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_135
timestamp 1
transform 1 0 13524 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636968456
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_153
timestamp 1
transform 1 0 15180 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_161
timestamp 1
transform 1 0 15916 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_176
timestamp 1
transform 1 0 17296 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_23
timestamp 1
transform 1 0 3220 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_33
timestamp 1
transform 1 0 4140 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_40
timestamp 1
transform 1 0 4784 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_57
timestamp 1
transform 1 0 6348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_63
timestamp 1
transform 1 0 6900 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_71
timestamp 1
transform 1 0 7636 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_84
timestamp 1636968456
transform 1 0 8832 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_113
timestamp 1
transform 1 0 11500 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_121
timestamp 1
transform 1 0 12236 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_131
timestamp 1
transform 1 0 13156 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_139
timestamp 1
transform 1 0 13892 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_148
timestamp 1
transform 1 0 14720 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_157
timestamp 1
transform 1 0 15548 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_161
timestamp 1
transform 1 0 15916 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_172
timestamp 1
transform 1 0 16928 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_178
timestamp 1
transform 1 0 17480 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_6
timestamp 1636968456
transform 1 0 1656 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_18
timestamp 1
transform 1 0 2760 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_29
timestamp 1
transform 1 0 3772 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_33
timestamp 1
transform 1 0 4140 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_40
timestamp 1
transform 1 0 4784 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_61
timestamp 1
transform 1 0 6716 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_85
timestamp 1
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_105
timestamp 1
transform 1 0 10764 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_118
timestamp 1
transform 1 0 11960 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_173
timestamp 1
transform 1 0 17020 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_6
timestamp 1
transform 1 0 1656 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636968456
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_40
timestamp 1
transform 1 0 4784 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_48
timestamp 1
transform 1 0 5520 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_64
timestamp 1
transform 1 0 6992 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_72
timestamp 1
transform 1 0 7728 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_77
timestamp 1
transform 1 0 8188 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_88
timestamp 1
transform 1 0 9200 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_94
timestamp 1
transform 1 0 9752 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_99
timestamp 1636968456
transform 1 0 10212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_113
timestamp 1
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_123
timestamp 1
transform 1 0 12420 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_129
timestamp 1636968456
transform 1 0 12972 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_141
timestamp 1
transform 1 0 14076 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1636968456
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_169
timestamp 1
transform 1 0 16652 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_177
timestamp 1
transform 1 0 17388 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp 1
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_35
timestamp 1636968456
transform 1 0 4324 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_47
timestamp 1636968456
transform 1 0 5428 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_59
timestamp 1
transform 1 0 6532 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_74
timestamp 1
transform 1 0 7912 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_85
timestamp 1
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_91
timestamp 1636968456
transform 1 0 9476 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_103
timestamp 1
transform 1 0 10580 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_107
timestamp 1
transform 1 0 10948 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_122
timestamp 1
transform 1 0 12328 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_130
timestamp 1
transform 1 0 13064 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_135
timestamp 1
transform 1 0 13524 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_141
timestamp 1
transform 1 0 14076 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_155
timestamp 1
transform 1 0 15364 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_163
timestamp 1
transform 1 0 16100 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_6
timestamp 1
transform 1 0 1656 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_15
timestamp 1
transform 1 0 2484 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_23
timestamp 1
transform 1 0 3220 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_42
timestamp 1636968456
transform 1 0 4968 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636968456
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1636968456
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_81
timestamp 1
transform 1 0 8556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_100
timestamp 1
transform 1 0 10304 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_113
timestamp 1
transform 1 0 11500 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_119
timestamp 1
transform 1 0 12052 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_143
timestamp 1
transform 1 0 14260 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_158
timestamp 1
transform 1 0 15640 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_176
timestamp 1
transform 1 0 17296 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_23
timestamp 1
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1636968456
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_41
timestamp 1
transform 1 0 4876 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_49
timestamp 1
transform 1 0 5612 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_57
timestamp 1
transform 1 0 6348 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_78
timestamp 1
transform 1 0 8280 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_85
timestamp 1
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_102
timestamp 1
transform 1 0 10488 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_131
timestamp 1
transform 1 0 13156 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_150
timestamp 1
transform 1 0 14904 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_158
timestamp 1
transform 1 0 15640 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_176
timestamp 1
transform 1 0 17296 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_6
timestamp 1
transform 1 0 1656 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_10
timestamp 1
transform 1 0 2024 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_14
timestamp 1
transform 1 0 2392 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_18
timestamp 1
transform 1 0 2760 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_26
timestamp 1636968456
transform 1 0 3496 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_38
timestamp 1
transform 1 0 4600 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp 1
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1
transform 1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_61
timestamp 1
transform 1 0 6716 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_73
timestamp 1636968456
transform 1 0 7820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_85
timestamp 1
transform 1 0 8924 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_94
timestamp 1636968456
transform 1 0 9752 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_106
timestamp 1
transform 1 0 10856 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1636968456
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1636968456
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1636968456
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_169
timestamp 1
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_177
timestamp 1
transform 1 0 17388 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_23
timestamp 1
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_36
timestamp 1
transform 1 0 4416 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_41
timestamp 1
transform 1 0 4876 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_57
timestamp 1
transform 1 0 6348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_68
timestamp 1
transform 1 0 7360 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1636968456
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1636968456
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1636968456
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_121
timestamp 1
transform 1 0 12236 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_126
timestamp 1636968456
transform 1 0 12696 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_146
timestamp 1
transform 1 0 14536 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_155
timestamp 1
transform 1 0 15364 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_163
timestamp 1
transform 1 0 16100 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_177
timestamp 1
transform 1 0 17388 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_6
timestamp 1
transform 1 0 1656 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_12
timestamp 1
transform 1 0 2208 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_16
timestamp 1
transform 1 0 2576 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_22
timestamp 1
transform 1 0 3128 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_48
timestamp 1
transform 1 0 5520 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_77
timestamp 1
transform 1 0 8188 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_106
timestamp 1
transform 1 0 10856 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_126
timestamp 1
transform 1 0 12696 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_178
timestamp 1
transform 1 0 17480 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_23
timestamp 1
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_35
timestamp 1636968456
transform 1 0 4324 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_47
timestamp 1636968456
transform 1 0 5428 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_62
timestamp 1636968456
transform 1 0 6808 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_74
timestamp 1
transform 1 0 7912 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_85
timestamp 1
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_93
timestamp 1
transform 1 0 9660 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_107
timestamp 1636968456
transform 1 0 10948 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_119
timestamp 1
transform 1 0 12052 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_131
timestamp 1
transform 1 0 13156 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_145
timestamp 1
transform 1 0 14444 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_154
timestamp 1
transform 1 0 15272 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_162
timestamp 1
transform 1 0 16008 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_176
timestamp 1
transform 1 0 17296 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_6
timestamp 1636968456
transform 1 0 1656 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_18
timestamp 1636968456
transform 1 0 2760 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_30
timestamp 1636968456
transform 1 0 3864 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_42
timestamp 1636968456
transform 1 0 4968 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_80
timestamp 1
transform 1 0 8464 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_88
timestamp 1
transform 1 0 9200 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_118
timestamp 1636968456
transform 1 0 11960 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_130
timestamp 1636968456
transform 1 0 13064 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_142
timestamp 1
transform 1 0 14168 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_150
timestamp 1
transform 1 0 14904 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_155
timestamp 1636968456
transform 1 0 15364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_173
timestamp 1
transform 1 0 17020 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_36
timestamp 1
transform 1 0 4416 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_49
timestamp 1
transform 1 0 5612 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_57
timestamp 1
transform 1 0 6348 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_67
timestamp 1
transform 1 0 7268 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_75
timestamp 1
transform 1 0 8004 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_92
timestamp 1
transform 1 0 9568 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_98
timestamp 1
transform 1 0 10120 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_106
timestamp 1636968456
transform 1 0 10856 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_118
timestamp 1
transform 1 0 11960 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_130
timestamp 1
transform 1 0 13064 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_141
timestamp 1
transform 1 0 14076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_147
timestamp 1
transform 1 0 14628 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_161
timestamp 1
transform 1 0 15916 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_168
timestamp 1
transform 1 0 16560 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_176
timestamp 1
transform 1 0 17296 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1636968456
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_15
timestamp 1
transform 1 0 2484 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_23
timestamp 1
transform 1 0 3220 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_41
timestamp 1636968456
transform 1 0 4876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp 1
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_57
timestamp 1
transform 1 0 6348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_66
timestamp 1
transform 1 0 7176 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_74
timestamp 1
transform 1 0 7912 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_89
timestamp 1
transform 1 0 9292 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_97
timestamp 1
transform 1 0 10028 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_102
timestamp 1
transform 1 0 10488 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_119
timestamp 1
transform 1 0 12052 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_133
timestamp 1
transform 1 0 13340 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_164
timestamp 1
transform 1 0 16192 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_177
timestamp 1
transform 1 0 17388 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_6
timestamp 1
transform 1 0 1656 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_10
timestamp 1
transform 1 0 2024 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_14
timestamp 1
transform 1 0 2392 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_29
timestamp 1
transform 1 0 3772 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_40
timestamp 1636968456
transform 1 0 4784 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_71
timestamp 1636968456
transform 1 0 7636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1636968456
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1636968456
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1636968456
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1636968456
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1636968456
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1636968456
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_165
timestamp 1
transform 1 0 16284 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_174
timestamp 1
transform 1 0 17112 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_178
timestamp 1
transform 1 0 17480 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_23
timestamp 1
transform 1 0 3220 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_28
timestamp 1
transform 1 0 3680 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_36
timestamp 1
transform 1 0 4416 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_50
timestamp 1
transform 1 0 5704 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_81
timestamp 1
transform 1 0 8556 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_113
timestamp 1
transform 1 0 11500 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_117
timestamp 1
transform 1 0 11868 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_144
timestamp 1
transform 1 0 14352 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_158
timestamp 1
transform 1 0 15640 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_162
timestamp 1
transform 1 0 16008 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_177
timestamp 1
transform 1 0 17388 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_6
timestamp 1
transform 1 0 1656 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_15
timestamp 1
transform 1 0 2484 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1636968456
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_50
timestamp 1
transform 1 0 5704 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_60
timestamp 1
transform 1 0 6624 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_163
timestamp 1
transform 1 0 16100 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_173
timestamp 1
transform 1 0 17020 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_23
timestamp 1636968456
transform 1 0 3220 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_35
timestamp 1636968456
transform 1 0 4324 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_47
timestamp 1
transform 1 0 5428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_64
timestamp 1636968456
transform 1 0 6992 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_76
timestamp 1
transform 1 0 8096 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_84
timestamp 1
transform 1 0 8832 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_91
timestamp 1
transform 1 0 9476 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_106
timestamp 1
transform 1 0 10856 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_113
timestamp 1
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_136
timestamp 1
transform 1 0 13616 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_176
timestamp 1
transform 1 0 17296 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_6
timestamp 1
transform 1 0 1656 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_12
timestamp 1
transform 1 0 2208 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_16
timestamp 1636968456
transform 1 0 2576 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_43
timestamp 1
transform 1 0 5060 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_62
timestamp 1636968456
transform 1 0 6808 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_74
timestamp 1
transform 1 0 7912 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp 1
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_93
timestamp 1
transform 1 0 9660 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_99
timestamp 1
transform 1 0 10212 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_113
timestamp 1636968456
transform 1 0 11500 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_125
timestamp 1636968456
transform 1 0 12604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_137
timestamp 1
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1636968456
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_153
timestamp 1
transform 1 0 15180 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_157
timestamp 1
transform 1 0 15548 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_23
timestamp 1
transform 1 0 3220 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_31
timestamp 1
transform 1 0 3956 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_41
timestamp 1636968456
transform 1 0 4876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1
transform 1 0 6348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_66
timestamp 1
transform 1 0 7176 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_72
timestamp 1
transform 1 0 7728 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_77
timestamp 1
transform 1 0 8188 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_85
timestamp 1
transform 1 0 8924 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_93
timestamp 1
transform 1 0 9660 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_113
timestamp 1
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_117
timestamp 1
transform 1 0 11868 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_129
timestamp 1
transform 1 0 12972 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_137
timestamp 1
transform 1 0 13708 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_155
timestamp 1
transform 1 0 15364 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_165
timestamp 1
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_172
timestamp 1
transform 1 0 16928 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_178
timestamp 1
transform 1 0 17480 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_23
timestamp 1
transform 1 0 3220 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1636968456
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_53
timestamp 1
transform 1 0 5980 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_65
timestamp 1
transform 1 0 7084 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_74
timestamp 1
transform 1 0 7912 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_93
timestamp 1
transform 1 0 9660 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_115
timestamp 1
transform 1 0 11684 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_119
timestamp 1
transform 1 0 12052 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_141
timestamp 1
transform 1 0 14076 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_156
timestamp 1
transform 1 0 15456 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_6
timestamp 1
transform 1 0 1656 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_10
timestamp 1
transform 1 0 2024 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_14
timestamp 1
transform 1 0 2392 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_18
timestamp 1
transform 1 0 2760 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_39
timestamp 1
transform 1 0 4692 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_43
timestamp 1
transform 1 0 5060 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_70
timestamp 1636968456
transform 1 0 7544 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_85
timestamp 1636968456
transform 1 0 8924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_97
timestamp 1636968456
transform 1 0 10028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_109
timestamp 1
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_113
timestamp 1
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_153
timestamp 1
transform 1 0 15180 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_157
timestamp 1
transform 1 0 15548 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_174
timestamp 1
transform 1 0 17112 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_178
timestamp 1
transform 1 0 17480 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_6
timestamp 1636968456
transform 1 0 1656 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_18
timestamp 1
transform 1 0 2760 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_37
timestamp 1636968456
transform 1 0 4508 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_49
timestamp 1636968456
transform 1 0 5612 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_61
timestamp 1636968456
transform 1 0 6716 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_73
timestamp 1
transform 1 0 7820 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_81
timestamp 1
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_85
timestamp 1
transform 1 0 8924 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_89
timestamp 1
transform 1 0 9292 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_118
timestamp 1
transform 1 0 11960 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_126
timestamp 1
transform 1 0 12696 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_141
timestamp 1
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_149
timestamp 1
transform 1 0 14812 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_158
timestamp 1
transform 1 0 15640 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_6
timestamp 1
transform 1 0 1656 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_10
timestamp 1
transform 1 0 2024 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_14
timestamp 1636968456
transform 1 0 2392 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_46
timestamp 1
transform 1 0 5336 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_60
timestamp 1
transform 1 0 6624 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_67
timestamp 1
transform 1 0 7268 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_73
timestamp 1
transform 1 0 7820 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_97
timestamp 1
transform 1 0 10028 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_105
timestamp 1
transform 1 0 10764 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_113
timestamp 1
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_121
timestamp 1
transform 1 0 12236 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_126
timestamp 1
transform 1 0 12696 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_152
timestamp 1
transform 1 0 15088 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_156
timestamp 1
transform 1 0 15456 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_160
timestamp 1
transform 1 0 15824 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_169
timestamp 1
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_177
timestamp 1
transform 1 0 17388 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_32
timestamp 1
transform 1 0 4048 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_88
timestamp 1
transform 1 0 9200 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_28_144
timestamp 1
transform 1 0 14352 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_170
timestamp 1
transform 1 0 16744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_174
timestamp 1
transform 1 0 17112 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_178
timestamp 1
transform 1 0 17480 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_9
timestamp 1
transform 1 0 1932 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_16
timestamp 1
transform 1 0 2576 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_24
timestamp 1
transform 1 0 3312 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_29
timestamp 1
transform 1 0 3772 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_40
timestamp 1
transform 1 0 4784 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_48
timestamp 1
transform 1 0 5520 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_52
timestamp 1
transform 1 0 5888 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_83
timestamp 1
transform 1 0 8740 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_88
timestamp 1
transform 1 0 9200 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_96
timestamp 1
transform 1 0 9936 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_100
timestamp 1
transform 1 0 10304 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_113
timestamp 1
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_124
timestamp 1
transform 1 0 12512 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_132
timestamp 1
transform 1 0 13248 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_136
timestamp 1
transform 1 0 13616 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_141
timestamp 1
transform 1 0 14076 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_148
timestamp 1
transform 1 0 14720 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_156
timestamp 1
transform 1 0 15456 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_160
timestamp 1
transform 1 0 15824 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_172
timestamp 1
transform 1 0 16928 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1
transform -1 0 1656 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1
transform -1 0 2576 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1
transform -1 0 3680 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1
transform -1 0 4784 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1
transform -1 0 5888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1
transform -1 0 6256 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1
transform 1 0 8464 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1
transform -1 0 9200 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1
transform 1 0 10028 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1
transform -1 0 11408 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1
transform -1 0 12512 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1
transform 1 0 13340 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1
transform -1 0 14720 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1
transform 1 0 15548 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1
transform 1 0 16652 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1
transform 1 0 17296 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  input17
timestamp 1
transform 1 0 9476 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  output18
timestamp 1
transform -1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output19
timestamp 1
transform -1 0 1656 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output20
timestamp 1
transform -1 0 1656 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output21
timestamp 1
transform -1 0 1656 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output22
timestamp 1
transform -1 0 1656 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output23
timestamp 1
transform -1 0 1656 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output24
timestamp 1
transform -1 0 1932 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output25
timestamp 1
transform -1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output26
timestamp 1
transform -1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output27
timestamp 1
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output28
timestamp 1
transform -1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output29
timestamp 1
transform -1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output30
timestamp 1
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output31
timestamp 1
transform -1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output32
timestamp 1
transform -1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  output33
timestamp 1
transform -1 0 1656 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_30
timestamp 1
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1
transform -1 0 17848 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_31
timestamp 1
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1
transform -1 0 17848 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_32
timestamp 1
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1
transform -1 0 17848 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_33
timestamp 1
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1
transform -1 0 17848 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_34
timestamp 1
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1
transform -1 0 17848 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_35
timestamp 1
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1
transform -1 0 17848 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_36
timestamp 1
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1
transform -1 0 17848 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_37
timestamp 1
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1
transform -1 0 17848 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_38
timestamp 1
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1
transform -1 0 17848 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_39
timestamp 1
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1
transform -1 0 17848 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_40
timestamp 1
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1
transform -1 0 17848 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_41
timestamp 1
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1
transform -1 0 17848 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_42
timestamp 1
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1
transform -1 0 17848 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_43
timestamp 1
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1
transform -1 0 17848 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_44
timestamp 1
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1
transform -1 0 17848 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_45
timestamp 1
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1
transform -1 0 17848 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_46
timestamp 1
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1
transform -1 0 17848 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_47
timestamp 1
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1
transform -1 0 17848 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_48
timestamp 1
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1
transform -1 0 17848 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_49
timestamp 1
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1
transform -1 0 17848 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_50
timestamp 1
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1
transform -1 0 17848 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_51
timestamp 1
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1
transform -1 0 17848 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_52
timestamp 1
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1
transform -1 0 17848 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_53
timestamp 1
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1
transform -1 0 17848 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_54
timestamp 1
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1
transform -1 0 17848 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_55
timestamp 1
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1
transform -1 0 17848 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_56
timestamp 1
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1
transform -1 0 17848 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_57
timestamp 1
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1
transform -1 0 17848 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_58
timestamp 1
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1
transform -1 0 17848 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_59
timestamp 1
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1
transform -1 0 17848 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_60
timestamp 1
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_61
timestamp 1
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_62
timestamp 1
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_63
timestamp 1
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_64
timestamp 1
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_65
timestamp 1
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_66
timestamp 1
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_67
timestamp 1
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_68
timestamp 1
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_69
timestamp 1
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_70
timestamp 1
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_71
timestamp 1
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_72
timestamp 1
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_73
timestamp 1
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_74
timestamp 1
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_75
timestamp 1
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_76
timestamp 1
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_77
timestamp 1
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_78
timestamp 1
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_79
timestamp 1
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_80
timestamp 1
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_81
timestamp 1
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_82
timestamp 1
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_83
timestamp 1
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_84
timestamp 1
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_85
timestamp 1
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_86
timestamp 1
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_87
timestamp 1
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_88
timestamp 1
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_89
timestamp 1
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_90
timestamp 1
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_91
timestamp 1
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_92
timestamp 1
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_93
timestamp 1
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_94
timestamp 1
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_95
timestamp 1
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_96
timestamp 1
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_97
timestamp 1
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_98
timestamp 1
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_99
timestamp 1
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_100
timestamp 1
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_101
timestamp 1
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_102
timestamp 1
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_103
timestamp 1
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_104
timestamp 1
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_105
timestamp 1
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_106
timestamp 1
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_107
timestamp 1
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_108
timestamp 1
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_109
timestamp 1
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_110
timestamp 1
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_111
timestamp 1
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_112
timestamp 1
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_113
timestamp 1
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_114
timestamp 1
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_115
timestamp 1
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_116
timestamp 1
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_117
timestamp 1
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_118
timestamp 1
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_119
timestamp 1
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_120
timestamp 1
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_121
timestamp 1
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_122
timestamp 1
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_123
timestamp 1
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_124
timestamp 1
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_125
timestamp 1
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_126
timestamp 1
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_127
timestamp 1
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_128
timestamp 1
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_129
timestamp 1
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_130
timestamp 1
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_131
timestamp 1
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_132
timestamp 1
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_133
timestamp 1
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_134
timestamp 1
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_135
timestamp 1
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_136
timestamp 1
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_137
timestamp 1
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_138
timestamp 1
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_139
timestamp 1
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_140
timestamp 1
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_141
timestamp 1
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_142
timestamp 1
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_143
timestamp 1
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_144
timestamp 1
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_145
timestamp 1
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_146
timestamp 1
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_147
timestamp 1
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_148
timestamp 1
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_149
timestamp 1
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_150
timestamp 1
transform 1 0 3680 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_151
timestamp 1
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_152
timestamp 1
transform 1 0 8832 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_153
timestamp 1
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_154
timestamp 1
transform 1 0 13984 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_155
timestamp 1
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
<< labels >>
flabel metal2 s 1122 20301 1178 21101 0 FreeSans 224 90 0 0 A[0]
port 0 nsew signal input
flabel metal2 s 2226 20301 2282 21101 0 FreeSans 224 90 0 0 A[1]
port 1 nsew signal input
flabel metal2 s 3330 20301 3386 21101 0 FreeSans 224 90 0 0 A[2]
port 2 nsew signal input
flabel metal2 s 4434 20301 4490 21101 0 FreeSans 224 90 0 0 A[3]
port 3 nsew signal input
flabel metal2 s 5538 20301 5594 21101 0 FreeSans 224 90 0 0 A[4]
port 4 nsew signal input
flabel metal2 s 6642 20301 6698 21101 0 FreeSans 224 90 0 0 A[5]
port 5 nsew signal input
flabel metal2 s 7746 20301 7802 21101 0 FreeSans 224 90 0 0 A[6]
port 6 nsew signal input
flabel metal2 s 8850 20301 8906 21101 0 FreeSans 224 90 0 0 A[7]
port 7 nsew signal input
flabel metal2 s 9954 20301 10010 21101 0 FreeSans 224 90 0 0 B[0]
port 8 nsew signal input
flabel metal2 s 11058 20301 11114 21101 0 FreeSans 224 90 0 0 B[1]
port 9 nsew signal input
flabel metal2 s 12162 20301 12218 21101 0 FreeSans 224 90 0 0 B[2]
port 10 nsew signal input
flabel metal2 s 13266 20301 13322 21101 0 FreeSans 224 90 0 0 B[3]
port 11 nsew signal input
flabel metal2 s 14370 20301 14426 21101 0 FreeSans 224 90 0 0 B[4]
port 12 nsew signal input
flabel metal2 s 15474 20301 15530 21101 0 FreeSans 224 90 0 0 B[5]
port 13 nsew signal input
flabel metal2 s 16578 20301 16634 21101 0 FreeSans 224 90 0 0 B[6]
port 14 nsew signal input
flabel metal2 s 17682 20301 17738 21101 0 FreeSans 224 90 0 0 B[7]
port 15 nsew signal input
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 Output[0]
port 16 nsew signal output
flabel metal3 s 0 13064 800 13184 0 FreeSans 480 0 0 0 Output[10]
port 17 nsew signal output
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 Output[11]
port 18 nsew signal output
flabel metal3 s 0 15240 800 15360 0 FreeSans 480 0 0 0 Output[12]
port 19 nsew signal output
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 Output[13]
port 20 nsew signal output
flabel metal3 s 0 17416 800 17536 0 FreeSans 480 0 0 0 Output[14]
port 21 nsew signal output
flabel metal3 s 0 18504 800 18624 0 FreeSans 480 0 0 0 Output[15]
port 22 nsew signal output
flabel metal3 s 0 3272 800 3392 0 FreeSans 480 0 0 0 Output[1]
port 23 nsew signal output
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 Output[2]
port 24 nsew signal output
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 Output[3]
port 25 nsew signal output
flabel metal3 s 0 6536 800 6656 0 FreeSans 480 0 0 0 Output[4]
port 26 nsew signal output
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 Output[5]
port 27 nsew signal output
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 Output[6]
port 28 nsew signal output
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 Output[7]
port 29 nsew signal output
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 Output[8]
port 30 nsew signal output
flabel metal3 s 0 11976 800 12096 0 FreeSans 480 0 0 0 Output[9]
port 31 nsew signal output
flabel metal4 s 2644 2128 3044 18544 0 FreeSans 1920 90 0 0 VGND
port 32 nsew ground bidirectional
flabel metal4 s 8644 2128 9044 18544 0 FreeSans 1920 90 0 0 VGND
port 32 nsew ground bidirectional
flabel metal4 s 14644 2128 15044 18544 0 FreeSans 1920 90 0 0 VGND
port 32 nsew ground bidirectional
flabel metal5 s 1056 3716 17896 4116 0 FreeSans 2560 0 0 0 VGND
port 32 nsew ground bidirectional
flabel metal5 s 1056 9716 17896 10116 0 FreeSans 2560 0 0 0 VGND
port 32 nsew ground bidirectional
flabel metal5 s 1056 15716 17896 16116 0 FreeSans 2560 0 0 0 VGND
port 32 nsew ground bidirectional
flabel metal4 s 1904 2128 2304 18544 0 FreeSans 1920 90 0 0 VPWR
port 33 nsew power bidirectional
flabel metal4 s 7904 2128 8304 18544 0 FreeSans 1920 90 0 0 VPWR
port 33 nsew power bidirectional
flabel metal4 s 13904 2128 14304 18544 0 FreeSans 1920 90 0 0 VPWR
port 33 nsew power bidirectional
flabel metal5 s 1056 2976 17896 3376 0 FreeSans 2560 0 0 0 VPWR
port 33 nsew power bidirectional
flabel metal5 s 1056 8976 17896 9376 0 FreeSans 2560 0 0 0 VPWR
port 33 nsew power bidirectional
flabel metal5 s 1056 14976 17896 15376 0 FreeSans 2560 0 0 0 VPWR
port 33 nsew power bidirectional
flabel metal3 s 18157 10344 18957 10464 0 FreeSans 480 0 0 0 clk
port 34 nsew signal input
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 reset
port 35 nsew signal input
rlabel metal1 9476 18496 9476 18496 0 VGND
rlabel metal1 9476 17952 9476 17952 0 VPWR
rlabel metal1 1288 18258 1288 18258 0 A[0]
rlabel metal1 2300 18258 2300 18258 0 A[1]
rlabel metal1 3404 18258 3404 18258 0 A[2]
rlabel metal1 4508 18258 4508 18258 0 A[3]
rlabel metal1 5612 18258 5612 18258 0 A[4]
rlabel metal1 6026 18292 6026 18292 0 A[5]
rlabel metal1 8326 18258 8326 18258 0 A[6]
rlabel metal1 9062 18258 9062 18258 0 A[7]
rlabel metal2 16054 14841 16054 14841 0 A_ff\[0\]
rlabel metal1 15134 10030 15134 10030 0 A_ff\[1\]
rlabel metal1 13110 11696 13110 11696 0 A_ff\[2\]
rlabel metal2 12834 13090 12834 13090 0 A_ff\[3\]
rlabel metal1 12558 12852 12558 12852 0 A_ff\[4\]
rlabel metal1 13984 6766 13984 6766 0 A_ff\[5\]
rlabel metal2 8602 6426 8602 6426 0 A_ff\[6\]
rlabel metal2 13110 13362 13110 13362 0 A_ff\[7\]
rlabel metal2 3910 3230 3910 3230 0 Adder.cla_16_bit.Sum\[0\]
rlabel metal1 3358 12682 3358 12682 0 Adder.cla_16_bit.Sum\[10\]
rlabel metal1 2944 13498 2944 13498 0 Adder.cla_16_bit.Sum\[11\]
rlabel metal1 3450 14586 3450 14586 0 Adder.cla_16_bit.Sum\[12\]
rlabel metal1 2898 15368 2898 15368 0 Adder.cla_16_bit.Sum\[13\]
rlabel metal1 3910 16762 3910 16762 0 Adder.cla_16_bit.Sum\[14\]
rlabel metal1 4002 16422 4002 16422 0 Adder.cla_16_bit.Sum\[15\]
rlabel metal1 6256 2958 6256 2958 0 Adder.cla_16_bit.Sum\[1\]
rlabel metal1 5244 2346 5244 2346 0 Adder.cla_16_bit.Sum\[2\]
rlabel metal1 3726 4012 3726 4012 0 Adder.cla_16_bit.Sum\[3\]
rlabel metal1 3542 5100 3542 5100 0 Adder.cla_16_bit.Sum\[4\]
rlabel metal2 3634 6460 3634 6460 0 Adder.cla_16_bit.Sum\[5\]
rlabel metal2 3450 7548 3450 7548 0 Adder.cla_16_bit.Sum\[6\]
rlabel metal1 2990 8398 2990 8398 0 Adder.cla_16_bit.Sum\[7\]
rlabel metal1 3358 10098 3358 10098 0 Adder.cla_16_bit.Sum\[8\]
rlabel metal1 2990 11186 2990 11186 0 Adder.cla_16_bit.Sum\[9\]
rlabel metal1 10120 18258 10120 18258 0 B[0]
rlabel metal2 11178 18751 11178 18751 0 B[1]
rlabel metal1 12236 18258 12236 18258 0 B[2]
rlabel metal1 13432 18258 13432 18258 0 B[3]
rlabel metal1 14444 18258 14444 18258 0 B[4]
rlabel metal1 15640 18258 15640 18258 0 B[5]
rlabel metal1 16744 18258 16744 18258 0 B[6]
rlabel metal1 17618 18258 17618 18258 0 B[7]
rlabel metal1 11638 17578 11638 17578 0 B_ff\[0\]
rlabel metal2 7498 6222 7498 6222 0 B_ff\[1\]
rlabel metal2 13662 5678 13662 5678 0 B_ff\[2\]
rlabel metal1 16974 13906 16974 13906 0 B_ff\[3\]
rlabel metal1 17342 13702 17342 13702 0 B_ff\[4\]
rlabel metal1 16974 12750 16974 12750 0 B_ff\[5\]
rlabel metal2 15870 16252 15870 16252 0 B_ff\[6\]
rlabel metal1 15594 15470 15594 15470 0 B_ff\[7\]
rlabel metal3 1050 2244 1050 2244 0 Output[0]
rlabel metal3 751 13124 751 13124 0 Output[10]
rlabel metal3 751 14212 751 14212 0 Output[11]
rlabel metal3 751 15300 751 15300 0 Output[12]
rlabel metal3 751 16388 751 16388 0 Output[13]
rlabel metal1 1380 17306 1380 17306 0 Output[14]
rlabel metal1 1472 18394 1472 18394 0 Output[15]
rlabel metal3 751 3332 751 3332 0 Output[1]
rlabel metal3 751 4420 751 4420 0 Output[2]
rlabel metal3 1050 5508 1050 5508 0 Output[3]
rlabel metal1 1380 6426 1380 6426 0 Output[4]
rlabel metal1 1380 7514 1380 7514 0 Output[5]
rlabel metal1 1380 8602 1380 8602 0 Output[6]
rlabel metal1 1380 9418 1380 9418 0 Output[7]
rlabel metal1 1380 10778 1380 10778 0 Output[8]
rlabel metal3 751 12036 751 12036 0 Output[9]
rlabel metal1 3680 2618 3680 2618 0 _000_
rlabel metal1 5336 2618 5336 2618 0 _001_
rlabel metal1 2300 2822 2300 2822 0 _002_
rlabel metal1 2905 4182 2905 4182 0 _003_
rlabel metal2 2346 5032 2346 5032 0 _004_
rlabel metal2 2346 6562 2346 6562 0 _005_
rlabel metal2 2346 7650 2346 7650 0 _006_
rlabel metal2 2254 8738 2254 8738 0 _007_
rlabel metal2 2438 9792 2438 9792 0 _008_
rlabel metal1 2905 11050 2905 11050 0 _009_
rlabel metal1 2300 12410 2300 12410 0 _010_
rlabel metal2 2346 13736 2346 13736 0 _011_
rlabel metal2 2438 14824 2438 14824 0 _012_
rlabel metal2 2346 15640 2346 15640 0 _013_
rlabel metal2 3910 16830 3910 16830 0 _014_
rlabel metal2 4462 17374 4462 17374 0 _015_
rlabel metal2 2254 17442 2254 17442 0 _016_
rlabel metal2 6670 10472 6670 10472 0 _017_
rlabel metal2 6486 17442 6486 17442 0 _018_
rlabel metal2 7130 17816 7130 17816 0 _019_
rlabel metal1 8142 17721 8142 17721 0 _020_
rlabel metal1 12604 17306 12604 17306 0 _021_
rlabel metal1 9200 16762 9200 16762 0 _022_
rlabel metal1 11086 16966 11086 16966 0 _023_
rlabel metal2 11086 17816 11086 17816 0 _024_
rlabel metal2 12466 8058 12466 8058 0 _025_
rlabel metal1 13478 6834 13478 6834 0 _026_
rlabel metal1 14260 17510 14260 17510 0 _027_
rlabel metal1 16744 14790 16744 14790 0 _028_
rlabel metal2 15686 17442 15686 17442 0 _029_
rlabel metal2 17066 17000 17066 17000 0 _030_
rlabel metal1 16889 15402 16889 15402 0 _031_
rlabel metal1 12972 4998 12972 4998 0 _032_
rlabel metal2 12282 3910 12282 3910 0 _033_
rlabel metal1 7038 4012 7038 4012 0 _034_
rlabel metal2 6210 4284 6210 4284 0 _035_
rlabel metal1 6532 4182 6532 4182 0 _036_
rlabel metal2 6394 3740 6394 3740 0 _037_
rlabel metal2 5934 4624 5934 4624 0 _038_
rlabel metal2 4554 3842 4554 3842 0 _039_
rlabel metal1 4048 5202 4048 5202 0 _040_
rlabel metal1 15962 12818 15962 12818 0 _041_
rlabel metal1 16192 11526 16192 11526 0 _042_
rlabel metal2 13938 13056 13938 13056 0 _043_
rlabel via2 15594 12835 15594 12835 0 _044_
rlabel metal1 16882 11526 16882 11526 0 _045_
rlabel metal1 14766 13940 14766 13940 0 _046_
rlabel metal1 17020 9894 17020 9894 0 _047_
rlabel metal2 16974 10234 16974 10234 0 _048_
rlabel metal2 16698 8177 16698 8177 0 _049_
rlabel metal1 8648 4250 8648 4250 0 _050_
rlabel metal1 10166 4692 10166 4692 0 _051_
rlabel metal1 11178 3502 11178 3502 0 _052_
rlabel metal2 10626 3332 10626 3332 0 _053_
rlabel metal1 10626 4590 10626 4590 0 _054_
rlabel metal1 10810 4794 10810 4794 0 _055_
rlabel metal1 10304 5542 10304 5542 0 _056_
rlabel metal1 10710 5542 10710 5542 0 _057_
rlabel via1 9890 5814 9890 5814 0 _058_
rlabel metal1 10166 5882 10166 5882 0 _059_
rlabel metal2 6670 5304 6670 5304 0 _060_
rlabel metal2 5474 4998 5474 4998 0 _061_
rlabel metal1 4922 5202 4922 5202 0 _062_
rlabel via1 4645 5202 4645 5202 0 _063_
rlabel metal1 4186 5134 4186 5134 0 _064_
rlabel metal1 15134 11220 15134 11220 0 _065_
rlabel metal1 15594 13974 15594 13974 0 _066_
rlabel metal1 16652 9554 16652 9554 0 _067_
rlabel metal2 14766 13226 14766 13226 0 _068_
rlabel metal1 15180 10778 15180 10778 0 _069_
rlabel metal2 17066 9180 17066 9180 0 _070_
rlabel metal1 16284 5746 16284 5746 0 _071_
rlabel metal1 15778 5134 15778 5134 0 _072_
rlabel metal1 16008 4998 16008 4998 0 _073_
rlabel via1 16790 4590 16790 4590 0 _074_
rlabel via1 15485 3502 15485 3502 0 _075_
rlabel metal2 15134 3264 15134 3264 0 _076_
rlabel metal1 15916 4658 15916 4658 0 _077_
rlabel metal1 16698 4794 16698 4794 0 _078_
rlabel metal1 16376 5338 16376 5338 0 _079_
rlabel metal2 16698 5236 16698 5236 0 _080_
rlabel metal1 16652 6766 16652 6766 0 _081_
rlabel metal2 16514 6103 16514 6103 0 _082_
rlabel metal1 7314 6222 7314 6222 0 _083_
rlabel metal1 5382 7378 5382 7378 0 _084_
rlabel metal2 6394 5950 6394 5950 0 _085_
rlabel metal1 6072 5882 6072 5882 0 _086_
rlabel metal2 4370 6086 4370 6086 0 _087_
rlabel metal2 4278 6086 4278 6086 0 _088_
rlabel metal2 13938 16388 13938 16388 0 _089_
rlabel metal1 15134 16048 15134 16048 0 _090_
rlabel metal1 15226 15436 15226 15436 0 _091_
rlabel metal1 16100 14858 16100 14858 0 _092_
rlabel metal2 15594 9724 15594 9724 0 _093_
rlabel metal2 15042 9146 15042 9146 0 _094_
rlabel metal1 15226 7412 15226 7412 0 _095_
rlabel metal1 13662 6766 13662 6766 0 _096_
rlabel metal1 14490 7378 14490 7378 0 _097_
rlabel metal1 14122 3706 14122 3706 0 _098_
rlabel metal2 14858 3978 14858 3978 0 _099_
rlabel metal1 15134 6698 15134 6698 0 _100_
rlabel metal1 14858 6630 14858 6630 0 _101_
rlabel metal2 14582 7242 14582 7242 0 _102_
rlabel metal1 15042 7310 15042 7310 0 _103_
rlabel metal2 15778 7684 15778 7684 0 _104_
rlabel metal1 16514 7888 16514 7888 0 _105_
rlabel metal1 16192 7854 16192 7854 0 _106_
rlabel metal2 17250 7004 17250 7004 0 _107_
rlabel metal2 10166 8160 10166 8160 0 _108_
rlabel metal1 4784 7378 4784 7378 0 _109_
rlabel metal1 4416 6766 4416 6766 0 _110_
rlabel metal1 4094 7344 4094 7344 0 _111_
rlabel metal2 3818 6596 3818 6596 0 _112_
rlabel metal1 3818 9112 3818 9112 0 _113_
rlabel metal1 13294 9452 13294 9452 0 _114_
rlabel metal2 12742 15164 12742 15164 0 _115_
rlabel metal1 12696 8942 12696 8942 0 _116_
rlabel metal2 12650 9350 12650 9350 0 _117_
rlabel metal2 15134 15538 15134 15538 0 _118_
rlabel metal1 13754 16048 13754 16048 0 _119_
rlabel metal1 12282 9452 12282 9452 0 _120_
rlabel metal1 12466 15028 12466 15028 0 _121_
rlabel metal1 13892 16150 13892 16150 0 _122_
rlabel metal1 11914 9554 11914 9554 0 _123_
rlabel metal2 12558 9724 12558 9724 0 _124_
rlabel metal1 6348 8942 6348 8942 0 _125_
rlabel via2 14398 6851 14398 6851 0 _126_
rlabel metal2 9798 7106 9798 7106 0 _127_
rlabel metal1 10672 7378 10672 7378 0 _128_
rlabel metal2 10166 7650 10166 7650 0 _129_
rlabel metal2 12650 5780 12650 5780 0 _130_
rlabel metal1 12742 5712 12742 5712 0 _131_
rlabel metal2 9982 7174 9982 7174 0 _132_
rlabel metal2 9614 7990 9614 7990 0 _133_
rlabel metal2 9982 8228 9982 8228 0 _134_
rlabel metal2 9522 7684 9522 7684 0 _135_
rlabel via2 15778 9571 15778 9571 0 _136_
rlabel metal1 15042 9146 15042 9146 0 _137_
rlabel metal1 14536 10166 14536 10166 0 _138_
rlabel metal2 13386 9248 13386 9248 0 _139_
rlabel metal1 7774 7752 7774 7752 0 _140_
rlabel metal1 7774 7990 7774 7990 0 _141_
rlabel metal1 7406 8058 7406 8058 0 _142_
rlabel metal2 7222 8228 7222 8228 0 _143_
rlabel metal1 7774 8500 7774 8500 0 _144_
rlabel metal1 6394 8466 6394 8466 0 _145_
rlabel metal1 5106 8942 5106 8942 0 _146_
rlabel metal2 5566 8466 5566 8466 0 _147_
rlabel metal2 5290 8976 5290 8976 0 _148_
rlabel metal2 4002 8602 4002 8602 0 _149_
rlabel metal2 12926 9724 12926 9724 0 _150_
rlabel metal1 13708 9486 13708 9486 0 _151_
rlabel metal1 9476 9554 9476 9554 0 _152_
rlabel metal1 15502 11084 15502 11084 0 _153_
rlabel metal1 14352 11118 14352 11118 0 _154_
rlabel metal1 12926 11016 12926 11016 0 _155_
rlabel metal1 11316 13362 11316 13362 0 _156_
rlabel metal2 14306 5508 14306 5508 0 _157_
rlabel metal2 14398 5644 14398 5644 0 _158_
rlabel metal1 11914 10608 11914 10608 0 _159_
rlabel metal1 10534 10064 10534 10064 0 _160_
rlabel metal2 10902 10234 10902 10234 0 _161_
rlabel metal1 10166 9656 10166 9656 0 _162_
rlabel metal1 9522 9418 9522 9418 0 _163_
rlabel metal2 9246 8976 9246 8976 0 _164_
rlabel metal1 8372 9146 8372 9146 0 _165_
rlabel metal2 8694 9146 8694 9146 0 _166_
rlabel metal1 7038 11084 7038 11084 0 _167_
rlabel metal2 7314 9146 7314 9146 0 _168_
rlabel metal1 7130 8908 7130 8908 0 _169_
rlabel metal1 5382 11084 5382 11084 0 _170_
rlabel metal1 4554 8976 4554 8976 0 _171_
rlabel metal1 4186 9554 4186 9554 0 _172_
rlabel metal1 4370 9588 4370 9588 0 _173_
rlabel metal1 4094 8942 4094 8942 0 _174_
rlabel metal1 4324 9146 4324 9146 0 _175_
rlabel metal1 3588 9690 3588 9690 0 _176_
rlabel metal1 13018 11764 13018 11764 0 _177_
rlabel metal2 13018 11356 13018 11356 0 _178_
rlabel metal1 9338 11084 9338 11084 0 _179_
rlabel metal2 9798 10948 9798 10948 0 _180_
rlabel metal1 12742 5236 12742 5236 0 _181_
rlabel metal2 12834 5644 12834 5644 0 _182_
rlabel metal1 11822 11526 11822 11526 0 _183_
rlabel metal2 10810 11526 10810 11526 0 _184_
rlabel metal1 14536 11866 14536 11866 0 _185_
rlabel metal1 14948 11730 14948 11730 0 _186_
rlabel metal1 11730 11662 11730 11662 0 _187_
rlabel metal1 9108 11730 9108 11730 0 _188_
rlabel metal1 9016 11186 9016 11186 0 _189_
rlabel metal1 8234 11764 8234 11764 0 _190_
rlabel metal2 7590 12002 7590 12002 0 _191_
rlabel metal1 7130 11220 7130 11220 0 _192_
rlabel metal2 6210 12036 6210 12036 0 _193_
rlabel metal1 6118 11118 6118 11118 0 _194_
rlabel metal2 5520 12818 5520 12818 0 _195_
rlabel metal2 4830 11526 4830 11526 0 _196_
rlabel metal2 4554 11968 4554 11968 0 _197_
rlabel metal1 4002 11186 4002 11186 0 _198_
rlabel metal2 4186 11968 4186 11968 0 _199_
rlabel metal2 11362 13532 11362 13532 0 _200_
rlabel metal2 11178 13940 11178 13940 0 _201_
rlabel metal1 14766 12920 14766 12920 0 _202_
rlabel metal1 15180 12886 15180 12886 0 _203_
rlabel metal1 16008 11866 16008 11866 0 _204_
rlabel metal2 11270 13260 11270 13260 0 _205_
rlabel metal1 10580 13974 10580 13974 0 _206_
rlabel metal2 11086 14688 11086 14688 0 _207_
rlabel metal2 10718 13260 10718 13260 0 _208_
rlabel metal1 9479 13838 9479 13838 0 _209_
rlabel metal1 10856 11798 10856 11798 0 _210_
rlabel metal1 8234 12784 8234 12784 0 _211_
rlabel metal1 8188 13294 8188 13294 0 _212_
rlabel metal1 12282 12852 12282 12852 0 _213_
rlabel metal1 13294 12750 13294 12750 0 _214_
rlabel metal1 9338 13906 9338 13906 0 _215_
rlabel metal1 7866 13498 7866 13498 0 _216_
rlabel metal1 6854 13294 6854 13294 0 _217_
rlabel metal1 6440 12206 6440 12206 0 _218_
rlabel metal1 4922 12750 4922 12750 0 _219_
rlabel metal1 4201 12818 4201 12818 0 _220_
rlabel metal1 4416 12682 4416 12682 0 _221_
rlabel metal1 3312 12410 3312 12410 0 _222_
rlabel metal1 3864 11730 3864 11730 0 _223_
rlabel metal2 3542 13124 3542 13124 0 _224_
rlabel metal2 8510 13260 8510 13260 0 _225_
rlabel metal1 6854 13906 6854 13906 0 _226_
rlabel metal2 14306 13090 14306 13090 0 _227_
rlabel metal2 15410 13498 15410 13498 0 _228_
rlabel metal1 15778 13328 15778 13328 0 _229_
rlabel metal1 14030 13430 14030 13430 0 _230_
rlabel metal2 9798 14212 9798 14212 0 _231_
rlabel metal2 10902 14756 10902 14756 0 _232_
rlabel metal2 10442 15232 10442 15232 0 _233_
rlabel metal1 10718 15436 10718 15436 0 _234_
rlabel metal1 10166 15028 10166 15028 0 _235_
rlabel metal2 12834 16252 12834 16252 0 _236_
rlabel metal2 12190 15436 12190 15436 0 _237_
rlabel metal1 10258 14892 10258 14892 0 _238_
rlabel metal1 7774 14382 7774 14382 0 _239_
rlabel metal1 6348 14382 6348 14382 0 _240_
rlabel metal2 6394 13498 6394 13498 0 _241_
rlabel metal1 5980 13498 5980 13498 0 _242_
rlabel metal1 5382 13396 5382 13396 0 _243_
rlabel metal1 4140 13362 4140 13362 0 _244_
rlabel metal1 14996 14994 14996 14994 0 _245_
rlabel metal1 14168 14994 14168 14994 0 _246_
rlabel metal1 11454 15504 11454 15504 0 _247_
rlabel metal2 11638 14756 11638 14756 0 _248_
rlabel metal1 10534 15674 10534 15674 0 _249_
rlabel metal1 9244 15470 9244 15470 0 _250_
rlabel metal2 8694 14688 8694 14688 0 _251_
rlabel metal1 7682 15538 7682 15538 0 _252_
rlabel metal1 8011 15470 8011 15470 0 _253_
rlabel metal1 6854 15368 6854 15368 0 _254_
rlabel metal1 7360 15062 7360 15062 0 _255_
rlabel metal2 6118 14586 6118 14586 0 _256_
rlabel metal2 5382 14654 5382 14654 0 _257_
rlabel metal1 5566 14348 5566 14348 0 _258_
rlabel metal1 5106 14314 5106 14314 0 _259_
rlabel metal1 4876 12274 4876 12274 0 _260_
rlabel metal1 4416 14586 4416 14586 0 _261_
rlabel metal2 5014 13770 5014 13770 0 _262_
rlabel metal2 4186 14314 4186 14314 0 _263_
rlabel metal1 4002 14416 4002 14416 0 _264_
rlabel metal1 13064 15130 13064 15130 0 _265_
rlabel metal1 12972 15470 12972 15470 0 _266_
rlabel metal2 9614 15674 9614 15674 0 _267_
rlabel metal1 7866 15028 7866 15028 0 _268_
rlabel metal2 7314 16150 7314 16150 0 _269_
rlabel metal1 8234 14994 8234 14994 0 _270_
rlabel metal2 7038 15130 7038 15130 0 _271_
rlabel metal1 5520 15470 5520 15470 0 _272_
rlabel viali 4737 15470 4737 15470 0 _273_
rlabel metal1 4324 15470 4324 15470 0 _274_
rlabel metal2 4278 15334 4278 15334 0 _275_
rlabel metal1 12673 15946 12673 15946 0 _276_
rlabel metal1 6808 16014 6808 16014 0 _277_
rlabel metal2 6578 16252 6578 16252 0 _278_
rlabel metal1 6210 16082 6210 16082 0 _279_
rlabel metal2 5842 16422 5842 16422 0 _280_
rlabel metal2 4094 16388 4094 16388 0 _281_
rlabel metal1 3266 16626 3266 16626 0 _282_
rlabel metal1 13202 4114 13202 4114 0 _283_
rlabel metal1 14674 9894 14674 9894 0 _284_
rlabel metal2 13478 15232 13478 15232 0 _285_
rlabel metal1 14352 14042 14352 14042 0 _286_
rlabel metal1 13846 13838 13846 13838 0 _287_
rlabel metal1 8034 3434 8034 3434 0 _288_
rlabel metal1 7360 2958 7360 2958 0 _289_
rlabel metal1 11868 6698 11868 6698 0 _290_
rlabel metal1 9016 4998 9016 4998 0 _291_
rlabel metal2 13846 5610 13846 5610 0 _292_
rlabel metal2 11546 6460 11546 6460 0 _293_
rlabel metal2 7682 6120 7682 6120 0 _294_
rlabel metal2 7912 5678 7912 5678 0 _295_
rlabel metal1 8372 3502 8372 3502 0 _296_
rlabel metal2 8326 3400 8326 3400 0 _297_
rlabel metal2 13754 3808 13754 3808 0 _298_
rlabel metal1 11316 2414 11316 2414 0 _299_
rlabel metal1 10396 2618 10396 2618 0 _300_
rlabel metal1 8786 2958 8786 2958 0 _301_
rlabel metal1 5428 4046 5428 4046 0 _302_
rlabel metal1 10718 2890 10718 2890 0 _303_
rlabel metal1 9656 3162 9656 3162 0 _304_
rlabel metal1 14904 5610 14904 5610 0 _305_
rlabel metal1 9154 3468 9154 3468 0 _306_
rlabel metal1 6302 3434 6302 3434 0 _307_
rlabel metal1 7682 5270 7682 5270 0 _308_
rlabel metal2 7222 4590 7222 4590 0 _309_
rlabel via1 12466 4114 12466 4114 0 _310_
rlabel metal1 13570 5780 13570 5780 0 _311_
rlabel metal2 11730 3366 11730 3366 0 _312_
rlabel metal2 16606 10557 16606 10557 0 clk
rlabel metal1 9292 12886 9292 12886 0 clknet_0_clk
rlabel metal1 3496 2482 3496 2482 0 clknet_2_0__leaf_clk
rlabel metal1 4922 12614 4922 12614 0 clknet_2_1__leaf_clk
rlabel metal1 5750 12750 5750 12750 0 clknet_2_2__leaf_clk
rlabel metal1 14628 14382 14628 14382 0 clknet_2_3__leaf_clk
rlabel metal1 1656 17578 1656 17578 0 net1
rlabel metal1 11592 18054 11592 18054 0 net10
rlabel metal3 12535 18020 12535 18020 0 net11
rlabel metal2 13294 17578 13294 17578 0 net12
rlabel metal1 15732 14314 15732 14314 0 net13
rlabel metal1 15272 17714 15272 17714 0 net14
rlabel metal2 16054 17340 16054 17340 0 net15
rlabel metal2 17250 16796 17250 16796 0 net16
rlabel metal1 4646 2414 4646 2414 0 net17
rlabel metal1 1610 2992 1610 2992 0 net18
rlabel metal2 1426 13124 1426 13124 0 net19
rlabel metal1 4140 18394 4140 18394 0 net2
rlabel metal2 1426 14212 1426 14212 0 net20
rlabel metal1 1518 15130 1518 15130 0 net21
rlabel metal2 1426 16116 1426 16116 0 net22
rlabel metal1 1610 17136 1610 17136 0 net23
rlabel metal1 1886 18224 1886 18224 0 net24
rlabel metal1 2185 3502 2185 3502 0 net25
rlabel metal1 1518 2618 1518 2618 0 net26
rlabel metal1 1472 4046 1472 4046 0 net27
rlabel metal1 1518 5338 1518 5338 0 net28
rlabel metal1 1518 6970 1518 6970 0 net29
rlabel metal2 4922 17816 4922 17816 0 net3
rlabel metal1 1518 8058 1518 8058 0 net30
rlabel metal2 1426 9350 1426 9350 0 net31
rlabel metal2 1426 10438 1426 10438 0 net32
rlabel metal2 1426 11764 1426 11764 0 net33
rlabel metal1 6578 18190 6578 18190 0 net4
rlabel metal2 7038 18054 7038 18054 0 net5
rlabel metal2 12190 17850 12190 17850 0 net6
rlabel metal1 8372 17238 8372 17238 0 net7
rlabel metal1 10064 16762 10064 16762 0 net8
rlabel metal2 10074 17884 10074 17884 0 net9
rlabel metal2 9430 1588 9430 1588 0 reset
<< properties >>
string FIXED_BBOX 0 0 18957 21101
<< end >>
